module leafVal1_rom
  #(
     parameter W_DATA = 11,
     parameter W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               8'b00000000: data1 <=  11'h216;
               8'b00000001: data1 <= -11'h1dd;
               8'b00000010: data1 <= -11'h182;
               8'b00000011: data1 <= -11'h0df;
               8'b00000100: data1 <= -11'h0c7;
               8'b00000101: data1 <=  11'h08e;
               8'b00000110: data1 <= -11'h1b0;
               8'b00000111: data1 <= -11'h17a;
               8'b00001000: data1 <= -11'h0db;
               8'b00001001: data1 <=  11'h13e;
               8'b00001010: data1 <= -11'h19e;
               8'b00001011: data1 <= -11'h1f1;
               8'b00001100: data1 <= -11'h08e;
               8'b00001101: data1 <=  11'h044;
               8'b00001110: data1 <= -11'h2ac;
               8'b00001111: data1 <= -11'h115;
               8'b00010000: data1 <= -11'h05a;
               8'b00010001: data1 <=  11'h0ed;
               8'b00010010: data1 <=  11'h128;
               8'b00010011: data1 <= -11'h06b;
               8'b00010100: data1 <=  11'h175;
               8'b00010101: data1 <=  11'h11e;
               8'b00010110: data1 <= -11'h059;
               8'b00010111: data1 <= -11'h09b;
               8'b00011000: data1 <=  11'h063;
               8'b00011001: data1 <= -11'h103;
               8'b00011010: data1 <= -11'h1a5;
               8'b00011011: data1 <=  11'h076;
               8'b00011100: data1 <= -11'h0a7;
               8'b00011101: data1 <= -11'h165;
               8'b00011110: data1 <= -11'h081;
               8'b00011111: data1 <=  11'h05d;
               8'b00100000: data1 <= -11'h04d;
               8'b00100001: data1 <= -11'h067;
               8'b00100010: data1 <=  11'h10d;
               8'b00100011: data1 <= -11'h1a0;
               8'b00100100: data1 <=  11'h048;
               8'b00100101: data1 <= -11'h103;
               8'b00100110: data1 <= -11'h02a;
               8'b00100111: data1 <=  11'h184;
               8'b00101000: data1 <=  11'h1c3;
               8'b00101001: data1 <= -11'h050;
               8'b00101010: data1 <= -11'h019;
               8'b00101011: data1 <= -11'h067;
               8'b00101100: data1 <=  11'h02b;
               8'b00101101: data1 <=  11'h0e3;
               8'b00101110: data1 <= -11'h05f;
               8'b00101111: data1 <=  11'h010;
               8'b00110000: data1 <= -11'h1bf;
               8'b00110001: data1 <= -11'h0f0;
               8'b00110010: data1 <= -11'h00d;
               8'b00110011: data1 <= -11'h1d4;
               8'b00110100: data1 <=  11'h127;
               8'b00110101: data1 <= -11'h190;
               8'b00110110: data1 <= -11'h093;
               8'b00110111: data1 <= -11'h175;
               8'b00111000: data1 <= -11'h0d5;
               8'b00111001: data1 <= -11'h050;
               8'b00111010: data1 <= -11'h06f;
               8'b00111011: data1 <=  11'h17d;
               8'b00111100: data1 <= -11'h0f6;
               8'b00111101: data1 <= -11'h272;
               8'b00111110: data1 <=  11'h02c;
               8'b00111111: data1 <=  11'h07c;
               8'b01000000: data1 <=  11'h02d;
               8'b01000001: data1 <= -11'h1f5;
               8'b01000010: data1 <=  11'h0fd;
               8'b01000011: data1 <= -11'h294;
               8'b01000100: data1 <=  11'h170;
               8'b01000101: data1 <= -11'h07e;
               8'b01000110: data1 <= -11'h254;
               8'b01000111: data1 <= -11'h0d8;
               8'b01001000: data1 <= -11'h171;
               8'b01001001: data1 <=  11'h02e;
               8'b01001010: data1 <=  11'h011;
               8'b01001011: data1 <=  11'h064;
               8'b01001100: data1 <=  11'h025;
               8'b01001101: data1 <=  11'h03f;
               8'b01001110: data1 <= -11'h0c1;
               8'b01001111: data1 <= -11'h05d;
               8'b01010000: data1 <= -11'h252;
               8'b01010001: data1 <=  11'h06c;
               8'b01010010: data1 <=  11'h11c;
               8'b01010011: data1 <= -11'h353;
               8'b01010100: data1 <= -11'h137;
               8'b01010101: data1 <= -11'h07b;
               8'b01010110: data1 <= -11'h114;
               8'b01010111: data1 <= -11'h133;
               8'b01011000: data1 <= -11'h070;
               8'b01011001: data1 <= -11'h02f;
               8'b01011010: data1 <=  11'h04d;
               8'b01011011: data1 <=  11'h13f;
               8'b01011100: data1 <= -11'h098;
               8'b01011101: data1 <=  11'h048;
               8'b01011110: data1 <=  11'h07b;
               8'b01011111: data1 <=  11'h044;
               8'b01100000: data1 <= -11'h14f;
               8'b01100001: data1 <=  11'h074;
               8'b01100010: data1 <= -11'h1bb;
               8'b01100011: data1 <= -11'h031;
               8'b01100100: data1 <= -11'h19c;
               8'b01100101: data1 <=  11'h0be;
               8'b01100110: data1 <= -11'h044;
               8'b01100111: data1 <= -11'h00f;
               8'b01101000: data1 <= -11'h059;
               8'b01101001: data1 <= -11'h10c;
               8'b01101010: data1 <=  11'h0d3;
               8'b01101011: data1 <=  11'h034;
               8'b01101100: data1 <=  11'h034;
               8'b01101101: data1 <= -11'h14c;
               8'b01101110: data1 <= -11'h14f;
               8'b01101111: data1 <= -11'h10d;
               8'b01110000: data1 <= -11'h15f;
               8'b01110001: data1 <= -11'h009;
               8'b01110010: data1 <= -11'h0ff;
               8'b01110011: data1 <=  11'h172;
               8'b01110100: data1 <= -11'h05f;
               8'b01110101: data1 <= -11'h093;
               8'b01110110: data1 <=  11'h004;
               8'b01110111: data1 <= -11'h014;
               8'b01111000: data1 <= -11'h126;
               8'b01111001: data1 <=  11'h05f;
               8'b01111010: data1 <=  11'h043;
               8'b01111011: data1 <=  11'h0c1;
               8'b01111100: data1 <=  11'h039;
               8'b01111101: data1 <= -11'h143;
               8'b01111110: data1 <=  11'h0de;
               8'b01111111: data1 <= -11'h163;
               8'b10000000: data1 <=  11'h010;
               8'b10000001: data1 <= -11'h089;
               8'b10000010: data1 <= -11'h05a;
               8'b10000011: data1 <= -11'h096;
               8'b10000100: data1 <= -11'h055;
               8'b10000101: data1 <=  11'h0b2;
               8'b10000110: data1 <=  11'h0dc;
               8'b10000111: data1 <=  11'h031;
               default: data1 <= 0;
           endcase
        end

endmodule: leafVal1_rom
