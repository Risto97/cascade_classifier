module leafVal0_rom
  #(
     W_DATA = 14,
     DEPTH = 2913,
     W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input ena,
     input [W_ADDR-1:0] addra,
     output [W_DATA-1:0] doa
    );

     (* rom_style = "block" *)


     logic [W_DATA-1:0] mem [DEPTH-1:0];

     always_ff @(posedge clk)
        begin
           if(ena)
              doa = mem[addra];
        end

     initial begin
         mem[0] = -14'h0237;
         mem[1] =  14'h0153;
         mem[2] =  14'h0110;
         mem[3] =  14'h012d;
         mem[4] =  14'h0142;
         mem[5] = -14'h01df;
         mem[6] =  14'h0070;
         mem[7] =  14'h0071;
         mem[8] =  14'h00da;
         mem[9] = -14'h0192;
         mem[10] =  14'h012e;
         mem[11] =  14'h00b3;
         mem[12] =  14'h01ba;
         mem[13] = -14'h022e;
         mem[14] =  14'h0074;
         mem[15] =  14'h0089;
         mem[16] =  14'h00ee;
         mem[17] = -14'h00a9;
         mem[18] = -14'h004c;
         mem[19] =  14'h015b;
         mem[20] = -14'h0032;
         mem[21] = -14'h0087;
         mem[22] =  14'h0124;
         mem[23] =  14'h00c5;
         mem[24] = -14'h0183;
         mem[25] =  14'h0177;
         mem[26] =  14'h0100;
         mem[27] = -14'h0198;
         mem[28] =  14'h00d4;
         mem[29] =  14'h006c;
         mem[30] =  14'h010d;
         mem[31] = -14'h0158;
         mem[32] =  14'h0173;
         mem[33] =  14'h0136;
         mem[34] = -14'h0075;
         mem[35] =  14'h0027;
         mem[36] = -14'h0190;
         mem[37] =  14'h003b;
         mem[38] =  14'h0147;
         mem[39] = -14'h004d;
         mem[40] = -14'h000d;
         mem[41] =  14'h0189;
         mem[42] =  14'h00ef;
         mem[43] =  14'h00f6;
         mem[44] = -14'h02f5;
         mem[45] = -14'h0070;
         mem[46] =  14'h0066;
         mem[47] = -14'h02a5;
         mem[48] =  14'h0048;
         mem[49] =  14'h003b;
         mem[50] =  14'h0113;
         mem[51] =  14'h0019;
         mem[52] = -14'h0112;
         mem[53] =  14'h00c4;
         mem[54] =  14'h0161;
         mem[55] =  14'h0084;
         mem[56] =  14'h0095;
         mem[57] =  14'h012b;
         mem[58] =  14'h00f4;
         mem[59] = -14'h0023;
         mem[60] =  14'h0046;
         mem[61] =  14'h003c;
         mem[62] = -14'h0157;
         mem[63] = -14'h00e6;
         mem[64] = -14'h01a2;
         mem[65] =  14'h002e;
         mem[66] = -14'h0061;
         mem[67] =  14'h003f;
         mem[68] = -14'h004b;
         mem[69] =  14'h00a1;
         mem[70] =  14'h000d;
         mem[71] =  14'h0063;
         mem[72] =  14'h0019;
         mem[73] = -14'h0142;
         mem[74] = -14'h0261;
         mem[75] = -14'h0046;
         mem[76] = -14'h0123;
         mem[77] = -14'h0144;
         mem[78] =  14'h0045;
         mem[79] =  14'h00b5;
         mem[80] =  14'h0009;
         mem[81] = -14'h000c;
         mem[82] = -14'h0059;
         mem[83] =  14'h0036;
         mem[84] =  14'h0115;
         mem[85] =  14'h0167;
         mem[86] =  14'h00bd;
         mem[87] =  14'h0060;
         mem[88] =  14'h0143;
         mem[89] =  14'h0075;
         mem[90] = -14'h00f5;
         mem[91] =  14'h000b;
         mem[92] =  14'h008a;
         mem[93] = -14'h017d;
         mem[94] = -14'h0086;
         mem[95] = -14'h0199;
         mem[96] =  14'h0027;
         mem[97] = -14'h00b8;
         mem[98] =  14'h0011;
         mem[99] =  14'h00ae;
         mem[100] =  14'h0013;
         mem[101] = -14'h0037;
         mem[102] =  14'h014f;
         mem[103] =  14'h0138;
         mem[104] =  14'h00d9;
         mem[105] =  14'h004c;
         mem[106] = -14'h0053;
         mem[107] = -14'h00d6;
         mem[108] = -14'h00ab;
         mem[109] =  14'h0023;
         mem[110] =  14'h0013;
         mem[111] =  14'h0031;
         mem[112] =  14'h0011;
         mem[113] =  14'h00c7;
         mem[114] =  14'h001f;
         mem[115] =  14'h0003;
         mem[116] =  14'h0087;
         mem[117] =  14'h0064;
         mem[118] = -14'h021e;
         mem[119] =  14'h00fc;
         mem[120] =  14'h0018;
         mem[121] = -14'h0025;
         mem[122] = -14'h0094;
         mem[123] = -14'h002b;
         mem[124] = -14'h00a3;
         mem[125] =  14'h0040;
         mem[126] = -14'h0045;
         mem[127] =  14'h003c;
         mem[128] = -14'h0143;
         mem[129] =  14'h004d;
         mem[130] =  14'h0087;
         mem[131] =  14'h003d;
         mem[132] =  14'h0084;
         mem[133] = -14'h0003;
         mem[134] = -14'h0042;
         mem[135] = -14'h0097;
         mem[136] =  14'h010b;
         mem[137] =  14'h008d;
         mem[138] =  14'h00a3;
         mem[139] =  14'h0088;
         mem[140] =  14'h005c;
         mem[141] =  14'h005c;
         mem[142] = -14'h0080;
         mem[143] =  14'h00da;
         mem[144] =  14'h0124;
         mem[145] = -14'h002e;
         mem[146] = -14'h0050;
         mem[147] =  14'h010b;
         mem[148] =  14'h0032;
         mem[149] = -14'h0154;
         mem[150] = -14'h00b3;
         mem[151] =  14'h0039;
         mem[152] = -14'h0083;
         mem[153] =  14'h009e;
         mem[154] =  14'h0079;
         mem[155] = -14'h00af;
         mem[156] =  14'h001d;
         mem[157] = -14'h000e;
         mem[158] =  14'h00d3;
         mem[159] = -14'h002d;
         mem[160] = -14'h018c;
         mem[161] =  14'h003d;
         mem[162] = -14'h0051;
         mem[163] = -14'h00d3;
         mem[164] =  14'h000d;
         mem[165] =  14'h0021;
         mem[166] =  14'h0009;
         mem[167] =  14'h007e;
         mem[168] = -14'h0092;
         mem[169] =  14'h00a3;
         mem[170] =  14'h0010;
         mem[171] = -14'h00ff;
         mem[172] =  14'h0009;
         mem[173] = -14'h010a;
         mem[174] = -14'h008a;
         mem[175] =  14'h0071;
         mem[176] =  14'h0000;
         mem[177] = -14'h00a5;
         mem[178] =  14'h00cd;
         mem[179] =  14'h0036;
         mem[180] = -14'h010e;
         mem[181] = -14'h00db;
         mem[182] =  14'h0010;
         mem[183] =  14'h00a2;
         mem[184] =  14'h0090;
         mem[185] = -14'h0181;
         mem[186] =  14'h0060;
         mem[187] =  14'h001f;
         mem[188] =  14'h00ad;
         mem[189] =  14'h00f3;
         mem[190] =  14'h007d;
         mem[191] =  14'h007f;
         mem[192] = -14'h0140;
         mem[193] =  14'h0098;
         mem[194] =  14'h004d;
         mem[195] =  14'h0039;
         mem[196] = -14'h0019;
         mem[197] =  14'h002f;
         mem[198] = -14'h0077;
         mem[199] = -14'h0043;
         mem[200] =  14'h006a;
         mem[201] =  14'h0097;
         mem[202] = -14'h0075;
         mem[203] =  14'h0024;
         mem[204] = -14'h00f9;
         mem[205] =  14'h002e;
         mem[206] = -14'h0153;
         mem[207] = -14'h0218;
         mem[208] =  14'h0083;
         mem[209] = -14'h0148;
         mem[210] = -14'h0076;
         mem[211] =  14'h000b;
         mem[212] =  14'h0058;
         mem[213] =  14'h006d;
         mem[214] =  14'h002a;
         mem[215] = -14'h0078;
         mem[216] = -14'h01ab;
         mem[217] =  14'h0009;
         mem[218] =  14'h003b;
         mem[219] =  14'h0019;
         mem[220] = -14'h0030;
         mem[221] = -14'h0061;
         mem[222] =  14'h0032;
         mem[223] =  14'h0081;
         mem[224] =  14'h003b;
         mem[225] = -14'h0051;
         mem[226] = -14'h0003;
         mem[227] =  14'h010a;
         mem[228] = -14'h00d5;
         mem[229] =  14'h0074;
         mem[230] = -14'h0180;
         mem[231] = -14'h0062;
         mem[232] = -14'h001b;
         mem[233] = -14'h01ae;
         mem[234] =  14'h003d;
         mem[235] =  14'h0077;
         mem[236] =  14'h002d;
         mem[237] =  14'h0012;
         mem[238] = -14'h018b;
         mem[239] =  14'h0060;
         mem[240] = -14'h013d;
         mem[241] =  14'h000d;
         mem[242] =  14'h003a;
         mem[243] =  14'h013a;
         mem[244] = -14'h000b;
         mem[245] = -14'h0037;
         mem[246] = -14'h01e6;
         mem[247] =  14'h0001;
         mem[248] = -14'h0015;
         mem[249] =  14'h0010;
         mem[250] = -14'h00c3;
         mem[251] =  14'h00d2;
         mem[252] =  14'h004b;
         mem[253] =  14'h0094;
         mem[254] =  14'h00e5;
         mem[255] =  14'h0081;
         mem[256] = -14'h00b4;
         mem[257] =  14'h00b5;
         mem[258] =  14'h0044;
         mem[259] = -14'h0062;
         mem[260] =  14'h0042;
         mem[261] = -14'h0096;
         mem[262] =  14'h002b;
         mem[263] = -14'h00e0;
         mem[264] =  14'h003c;
         mem[265] = -14'h0090;
         mem[266] =  14'h0062;
         mem[267] = -14'h0163;
         mem[268] = -14'h0111;
         mem[269] =  14'h0032;
         mem[270] =  14'h006f;
         mem[271] = -14'h0072;
         mem[272] =  14'h0039;
         mem[273] = -14'h0001;
         mem[274] = -14'h0085;
         mem[275] = -14'h0182;
         mem[276] =  14'h002f;
         mem[277] =  14'h0000;
         mem[278] = -14'h0238;
         mem[279] =  14'h000f;
         mem[280] = -14'h012f;
         mem[281] =  14'h001f;
         mem[282] =  14'h00b5;
         mem[283] = -14'h010d;
         mem[284] =  14'h0031;
         mem[285] = -14'h0040;
         mem[286] = -14'h0036;
         mem[287] = -14'h0047;
         mem[288] =  14'h003e;
         mem[289] =  14'h000e;
         mem[290] =  14'h0032;
         mem[291] =  14'h010d;
         mem[292] = -14'h01b8;
         mem[293] =  14'h000f;
         mem[294] =  14'h0007;
         mem[295] = -14'h007b;
         mem[296] =  14'h0029;
         mem[297] =  14'h000a;
         mem[298] =  14'h0052;
         mem[299] = -14'h0043;
         mem[300] =  14'h0026;
         mem[301] =  14'h000a;
         mem[302] =  14'h0027;
         mem[303] = -14'h006c;
         mem[304] =  14'h002f;
         mem[305] =  14'h0000;
         mem[306] =  14'h004f;
         mem[307] = -14'h00a6;
         mem[308] =  14'h0027;
         mem[309] =  14'h0187;
         mem[310] =  14'h00a6;
         mem[311] =  14'h0009;
         mem[312] = -14'h0019;
         mem[313] = -14'h0057;
         mem[314] = -14'h0004;
         mem[315] = -14'h0007;
         mem[316] =  14'h002a;
         mem[317] =  14'h0000;
         mem[318] = -14'h002d;
         mem[319] = -14'h0147;
         mem[320] = -14'h0184;
         mem[321] =  14'h0053;
         mem[322] =  14'h0026;
         mem[323] =  14'h011c;
         mem[324] = -14'h009d;
         mem[325] =  14'h0065;
         mem[326] =  14'h0049;
         mem[327] =  14'h0073;
         mem[328] = -14'h00ae;
         mem[329] =  14'h000f;
         mem[330] = -14'h01ba;
         mem[331] =  14'h001f;
         mem[332] = -14'h00cf;
         mem[333] =  14'h00ac;
         mem[334] =  14'h00d7;
         mem[335] = -14'h0079;
         mem[336] =  14'h00f2;
         mem[337] = -14'h0050;
         mem[338] =  14'h002d;
         mem[339] =  14'h003f;
         mem[340] = -14'h006d;
         mem[341] = -14'h0199;
         mem[342] =  14'h0060;
         mem[343] =  14'h003f;
         mem[344] = -14'h0171;
         mem[345] = -14'h015c;
         mem[346] =  14'h0045;
         mem[347] = -14'h00d0;
         mem[348] = -14'h00bf;
         mem[349] =  14'h00cf;
         mem[350] =  14'h00dc;
         mem[351] = -14'h00fd;
         mem[352] =  14'h0027;
         mem[353] = -14'h00b4;
         mem[354] = -14'h0067;
         mem[355] =  14'h0012;
         mem[356] = -14'h00b8;
         mem[357] =  14'h0043;
         mem[358] =  14'h0025;
         mem[359] = -14'h0113;
         mem[360] =  14'h0137;
         mem[361] =  14'h0003;
         mem[362] = -14'h0027;
         mem[363] =  14'h00b4;
         mem[364] =  14'h0055;
         mem[365] =  14'h0013;
         mem[366] =  14'h000c;
         mem[367] = -14'h003e;
         mem[368] =  14'h001f;
         mem[369] = -14'h0006;
         mem[370] = -14'h001e;
         mem[371] = -14'h0044;
         mem[372] = -14'h00a5;
         mem[373] = -14'h013d;
         mem[374] =  14'h0104;
         mem[375] = -14'h005c;
         mem[376] =  14'h0034;
         mem[377] = -14'h0005;
         mem[378] = -14'h004b;
         mem[379] =  14'h0115;
         mem[380] =  14'h0137;
         mem[381] = -14'h0110;
         mem[382] =  14'h002b;
         mem[383] =  14'h0084;
         mem[384] =  14'h003f;
         mem[385] = -14'h0250;
         mem[386] = -14'h0053;
         mem[387] =  14'h0012;
         mem[388] = -14'h01b9;
         mem[389] =  14'h0104;
         mem[390] =  14'h0026;
         mem[391] = -14'h004a;
         mem[392] = -14'h0056;
         mem[393] = -14'h0258;
         mem[394] =  14'h0027;
         mem[395] = -14'h0007;
         mem[396] =  14'h003c;
         mem[397] =  14'h00ec;
         mem[398] =  14'h004f;
         mem[399] = -14'h02b5;
         mem[400] = -14'h0008;
         mem[401] =  14'h003a;
         mem[402] = -14'h010b;
         mem[403] =  14'h00c4;
         mem[404] =  14'h0047;
         mem[405] = -14'h0041;
         mem[406] =  14'h0118;
         mem[407] =  14'h0087;
         mem[408] =  14'h0067;
         mem[409] =  14'h00bd;
         mem[410] =  14'h00bc;
         mem[411] =  14'h0061;
         mem[412] =  14'h005d;
         mem[413] =  14'h00cb;
         mem[414] = -14'h0054;
         mem[415] = -14'h00f7;
         mem[416] = -14'h010f;
         mem[417] =  14'h0022;
         mem[418] =  14'h009a;
         mem[419] = -14'h0036;
         mem[420] = -14'h0177;
         mem[421] =  14'h0034;
         mem[422] =  14'h001a;
         mem[423] = -14'h0066;
         mem[424] = -14'h019b;
         mem[425] = -14'h0022;
         mem[426] =  14'h0002;
         mem[427] =  14'h0042;
         mem[428] = -14'h00b7;
         mem[429] = -14'h01a5;
         mem[430] =  14'h0006;
         mem[431] = -14'h001a;
         mem[432] = -14'h0089;
         mem[433] =  14'h0033;
         mem[434] = -14'h0102;
         mem[435] = -14'h0046;
         mem[436] = -14'h0088;
         mem[437] =  14'h0035;
         mem[438] = -14'h0009;
         mem[439] = -14'h00b6;
         mem[440] =  14'h0004;
         mem[441] = -14'h0010;
         mem[442] =  14'h00cb;
         mem[443] = -14'h00af;
         mem[444] = -14'h0037;
         mem[445] =  14'h013f;
         mem[446] =  14'h0025;
         mem[447] = -14'h0003;
         mem[448] =  14'h0114;
         mem[449] =  14'h0123;
         mem[450] = -14'h0001;
         mem[451] =  14'h003d;
         mem[452] = -14'h0034;
         mem[453] = -14'h0138;
         mem[454] =  14'h000d;
         mem[455] =  14'h004a;
         mem[456] = -14'h00ab;
         mem[457] =  14'h0004;
         mem[458] =  14'h0006;
         mem[459] =  14'h0007;
         mem[460] =  14'h0097;
         mem[461] =  14'h0043;
         mem[462] = -14'h0055;
         mem[463] =  14'h0028;
         mem[464] = -14'h0006;
         mem[465] = -14'h000b;
         mem[466] = -14'h0072;
         mem[467] =  14'h0024;
         mem[468] = -14'h0061;
         mem[469] =  14'h0010;
         mem[470] =  14'h00cb;
         mem[471] =  14'h001d;
         mem[472] = -14'h0001;
         mem[473] =  14'h0068;
         mem[474] = -14'h0062;
         mem[475] =  14'h00c4;
         mem[476] = -14'h0039;
         mem[477] = -14'h0174;
         mem[478] =  14'h0042;
         mem[479] =  14'h007c;
         mem[480] = -14'h0038;
         mem[481] =  14'h0025;
         mem[482] = -14'h0033;
         mem[483] =  14'h0045;
         mem[484] = -14'h0030;
         mem[485] =  14'h0028;
         mem[486] = -14'h01a3;
         mem[487] =  14'h003d;
         mem[488] = -14'h0001;
         mem[489] = -14'h0073;
         mem[490] =  14'h0070;
         mem[491] =  14'h0040;
         mem[492] =  14'h0006;
         mem[493] =  14'h0000;
         mem[494] =  14'h0185;
         mem[495] = -14'h0037;
         mem[496] =  14'h0005;
         mem[497] =  14'h00a4;
         mem[498] =  14'h0093;
         mem[499] =  14'h0150;
         mem[500] =  14'h004a;
         mem[501] =  14'h0088;
         mem[502] = -14'h0072;
         mem[503] = -14'h0046;
         mem[504] =  14'h0034;
         mem[505] =  14'h0011;
         mem[506] = -14'h0085;
         mem[507] =  14'h000b;
         mem[508] =  14'h002f;
         mem[509] = -14'h00b0;
         mem[510] = -14'h00d7;
         mem[511] = -14'h015d;
         mem[512] =  14'h0042;
         mem[513] =  14'h0010;
         mem[514] = -14'h0004;
         mem[515] = -14'h0053;
         mem[516] =  14'h0033;
         mem[517] =  14'h0039;
         mem[518] = -14'h0112;
         mem[519] =  14'h0009;
         mem[520] = -14'h00b7;
         mem[521] = -14'h0088;
         mem[522] =  14'h00f9;
         mem[523] = -14'h003c;
         mem[524] =  14'h0075;
         mem[525] = -14'h02aa;
         mem[526] =  14'h0006;
         mem[527] = -14'h022b;
         mem[528] =  14'h00bf;
         mem[529] =  14'h0002;
         mem[530] =  14'h00fe;
         mem[531] = -14'h003f;
         mem[532] = -14'h009c;
         mem[533] =  14'h0007;
         mem[534] = -14'h0022;
         mem[535] = -14'h0085;
         mem[536] =  14'h0026;
         mem[537] =  14'h0000;
         mem[538] = -14'h009d;
         mem[539] = -14'h0035;
         mem[540] =  14'h007a;
         mem[541] =  14'h001c;
         mem[542] = -14'h017f;
         mem[543] =  14'h00d0;
         mem[544] = -14'h0011;
         mem[545] =  14'h000c;
         mem[546] = -14'h0001;
         mem[547] = -14'h002f;
         mem[548] =  14'h0018;
         mem[549] = -14'h0045;
         mem[550] =  14'h0028;
         mem[551] = -14'h003c;
         mem[552] =  14'h0032;
         mem[553] =  14'h0005;
         mem[554] = -14'h0004;
         mem[555] = -14'h01bc;
         mem[556] = -14'h000e;
         mem[557] = -14'h00c5;
         mem[558] =  14'h00ab;
         mem[559] =  14'h004f;
         mem[560] =  14'h0041;
         mem[561] =  14'h0069;
         mem[562] =  14'h0004;
         mem[563] = -14'h0035;
         mem[564] =  14'h000a;
         mem[565] =  14'h002b;
         mem[566] =  14'h00d1;
         mem[567] =  14'h0006;
         mem[568] = -14'h0057;
         mem[569] =  14'h0000;
         mem[570] =  14'h0040;
         mem[571] = -14'h016e;
         mem[572] =  14'h0055;
         mem[573] =  14'h0021;
         mem[574] = -14'h004f;
         mem[575] =  14'h00b5;
         mem[576] =  14'h0031;
         mem[577] = -14'h00e3;
         mem[578] = -14'h0046;
         mem[579] =  14'h0006;
         mem[580] = -14'h002c;
         mem[581] = -14'h0033;
         mem[582] =  14'h001d;
         mem[583] = -14'h0074;
         mem[584] =  14'h0064;
         mem[585] = -14'h0033;
         mem[586] =  14'h0034;
         mem[587] = -14'h0105;
         mem[588] = -14'h0017;
         mem[589] = -14'h01ed;
         mem[590] = -14'h0011;
         mem[591] =  14'h002f;
         mem[592] =  14'h0038;
         mem[593] = -14'h002f;
         mem[594] =  14'h005f;
         mem[595] = -14'h0044;
         mem[596] =  14'h0093;
         mem[597] =  14'h0102;
         mem[598] =  14'h0090;
         mem[599] =  14'h004f;
         mem[600] = -14'h011e;
         mem[601] =  14'h0054;
         mem[602] =  14'h0086;
         mem[603] = -14'h0008;
         mem[604] =  14'h001e;
         mem[605] =  14'h0035;
         mem[606] = -14'h0048;
         mem[607] = -14'h00b3;
         mem[608] =  14'h00bb;
         mem[609] =  14'h0027;
         mem[610] = -14'h0057;
         mem[611] = -14'h0021;
         mem[612] = -14'h00f5;
         mem[613] = -14'h0077;
         mem[614] = -14'h0086;
         mem[615] =  14'h0037;
         mem[616] =  14'h0010;
         mem[617] =  14'h0037;
         mem[618] =  14'h000c;
         mem[619] =  14'h002c;
         mem[620] = -14'h0038;
         mem[621] =  14'h002e;
         mem[622] =  14'h000e;
         mem[623] =  14'h0086;
         mem[624] =  14'h008f;
         mem[625] = -14'h00b3;
         mem[626] =  14'h000b;
         mem[627] =  14'h0042;
         mem[628] =  14'h0094;
         mem[629] =  14'h0032;
         mem[630] =  14'h0036;
         mem[631] =  14'h00c5;
         mem[632] = -14'h003f;
         mem[633] = -14'h0009;
         mem[634] =  14'h011a;
         mem[635] =  14'h00b8;
         mem[636] =  14'h000b;
         mem[637] = -14'h0060;
         mem[638] =  14'h011e;
         mem[639] =  14'h0031;
         mem[640] = -14'h0129;
         mem[641] =  14'h002a;
         mem[642] = -14'h0003;
         mem[643] = -14'h0015;
         mem[644] =  14'h0098;
         mem[645] =  14'h0022;
         mem[646] = -14'h0008;
         mem[647] =  14'h0004;
         mem[648] =  14'h0088;
         mem[649] =  14'h0029;
         mem[650] = -14'h00c0;
         mem[651] = -14'h00a7;
         mem[652] = -14'h013a;
         mem[653] =  14'h006e;
         mem[654] = -14'h0131;
         mem[655] =  14'h0024;
         mem[656] =  14'h008a;
         mem[657] =  14'h0090;
         mem[658] = -14'h00cb;
         mem[659] =  14'h017b;
         mem[660] = -14'h0007;
         mem[661] =  14'h0008;
         mem[662] =  14'h004c;
         mem[663] = -14'h0061;
         mem[664] = -14'h0087;
         mem[665] =  14'h021a;
         mem[666] = -14'h000a;
         mem[667] =  14'h005b;
         mem[668] = -14'h002d;
         mem[669] = -14'h014c;
         mem[670] =  14'h0023;
         mem[671] =  14'h0064;
         mem[672] = -14'h00b8;
         mem[673] =  14'h0010;
         mem[674] = -14'h002a;
         mem[675] = -14'h002a;
         mem[676] =  14'h00bb;
         mem[677] =  14'h0034;
         mem[678] = -14'h004b;
         mem[679] =  14'h0067;
         mem[680] = -14'h002c;
         mem[681] =  14'h00b2;
         mem[682] =  14'h0000;
         mem[683] =  14'h0089;
         mem[684] = -14'h00bf;
         mem[685] =  14'h0055;
         mem[686] = -14'h0009;
         mem[687] =  14'h0004;
         mem[688] =  14'h00ba;
         mem[689] = -14'h007d;
         mem[690] =  14'h00c5;
         mem[691] =  14'h0011;
         mem[692] = -14'h002f;
         mem[693] = -14'h019a;
         mem[694] =  14'h0130;
         mem[695] =  14'h0064;
         mem[696] = -14'h019c;
         mem[697] =  14'h008a;
         mem[698] = -14'h0051;
         mem[699] = -14'h0107;
         mem[700] = -14'h00ca;
         mem[701] = -14'h00d6;
         mem[702] = -14'h00a0;
         mem[703] =  14'h0192;
         mem[704] =  14'h0062;
         mem[705] =  14'h0086;
         mem[706] = -14'h0048;
         mem[707] = -14'h004e;
         mem[708] = -14'h00df;
         mem[709] = -14'h0033;
         mem[710] =  14'h0014;
         mem[711] =  14'h0091;
         mem[712] =  14'h0072;
         mem[713] =  14'h00ad;
         mem[714] =  14'h0031;
         mem[715] = -14'h00b6;
         mem[716] =  14'h001d;
         mem[717] =  14'h0033;
         mem[718] =  14'h005d;
         mem[719] =  14'h0020;
         mem[720] =  14'h0093;
         mem[721] = -14'h0086;
         mem[722] =  14'h007a;
         mem[723] = -14'h018e;
         mem[724] =  14'h0030;
         mem[725] = -14'h0072;
         mem[726] = -14'h0036;
         mem[727] =  14'h0085;
         mem[728] =  14'h0007;
         mem[729] = -14'h0039;
         mem[730] =  14'h0025;
         mem[731] =  14'h0004;
         mem[732] = -14'h00fc;
         mem[733] =  14'h0005;
         mem[734] =  14'h0032;
         mem[735] =  14'h0061;
         mem[736] = -14'h0025;
         mem[737] = -14'h0047;
         mem[738] =  14'h009a;
         mem[739] = -14'h0060;
         mem[740] =  14'h0108;
         mem[741] = -14'h0039;
         mem[742] = -14'h012f;
         mem[743] =  14'h000b;
         mem[744] =  14'h0112;
         mem[745] = -14'h002c;
         mem[746] = -14'h0012;
         mem[747] =  14'h0066;
         mem[748] = -14'h0137;
         mem[749] = -14'h00b6;
         mem[750] =  14'h002e;
         mem[751] = -14'h018b;
         mem[752] =  14'h002a;
         mem[753] = -14'h0004;
         mem[754] =  14'h003c;
         mem[755] =  14'h000e;
         mem[756] = -14'h0004;
         mem[757] = -14'h0036;
         mem[758] =  14'h002f;
         mem[759] = -14'h0065;
         mem[760] = -14'h0291;
         mem[761] = -14'h0003;
         mem[762] =  14'h002a;
         mem[763] =  14'h0054;
         mem[764] = -14'h007c;
         mem[765] = -14'h0039;
         mem[766] =  14'h0030;
         mem[767] = -14'h0035;
         mem[768] = -14'h0099;
         mem[769] = -14'h0005;
         mem[770] =  14'h000f;
         mem[771] = -14'h018a;
         mem[772] =  14'h005f;
         mem[773] =  14'h0023;
         mem[774] = -14'h0004;
         mem[775] = -14'h0139;
         mem[776] =  14'h0000;
         mem[777] = -14'h0003;
         mem[778] = -14'h013d;
         mem[779] =  14'h0083;
         mem[780] = -14'h00b5;
         mem[781] =  14'h0000;
         mem[782] =  14'h0025;
         mem[783] = -14'h0077;
         mem[784] = -14'h006a;
         mem[785] =  14'h006f;
         mem[786] = -14'h00f3;
         mem[787] = -14'h004e;
         mem[788] = -14'h01fa;
         mem[789] = -14'h0002;
         mem[790] = -14'h0008;
         mem[791] =  14'h0063;
         mem[792] =  14'h0096;
         mem[793] = -14'h00f2;
         mem[794] =  14'h0036;
         mem[795] = -14'h0007;
         mem[796] =  14'h0129;
         mem[797] = -14'h011d;
         mem[798] =  14'h0035;
         mem[799] = -14'h0028;
         mem[800] =  14'h002e;
         mem[801] =  14'h000b;
         mem[802] = -14'h00bf;
         mem[803] = -14'h01ac;
         mem[804] =  14'h00c3;
         mem[805] = -14'h00e2;
         mem[806] = -14'h0276;
         mem[807] = -14'h004c;
         mem[808] =  14'h0029;
         mem[809] = -14'h005f;
         mem[810] =  14'h0098;
         mem[811] =  14'h008d;
         mem[812] =  14'h0068;
         mem[813] = -14'h003c;
         mem[814] =  14'h0028;
         mem[815] = -14'h0057;
         mem[816] =  14'h0018;
         mem[817] =  14'h0008;
         mem[818] = -14'h000d;
         mem[819] = -14'h0005;
         mem[820] =  14'h00ea;
         mem[821] = -14'h0049;
         mem[822] =  14'h0088;
         mem[823] = -14'h0071;
         mem[824] = -14'h028f;
         mem[825] = -14'h011b;
         mem[826] =  14'h0091;
         mem[827] =  14'h0020;
         mem[828] =  14'h00df;
         mem[829] =  14'h0035;
         mem[830] =  14'h000e;
         mem[831] = -14'h0002;
         mem[832] =  14'h002b;
         mem[833] = -14'h0163;
         mem[834] =  14'h0000;
         mem[835] = -14'h006a;
         mem[836] =  14'h0004;
         mem[837] = -14'h0032;
         mem[838] =  14'h0084;
         mem[839] =  14'h00b4;
         mem[840] = -14'h00ab;
         mem[841] =  14'h005b;
         mem[842] =  14'h0030;
         mem[843] =  14'h0043;
         mem[844] =  14'h0044;
         mem[845] = -14'h0114;
         mem[846] = -14'h0047;
         mem[847] =  14'h003d;
         mem[848] = -14'h003f;
         mem[849] =  14'h0001;
         mem[850] =  14'h00b5;
         mem[851] = -14'h0170;
         mem[852] =  14'h000c;
         mem[853] = -14'h0072;
         mem[854] =  14'h0058;
         mem[855] = -14'h0157;
         mem[856] = -14'h0084;
         mem[857] = -14'h00ba;
         mem[858] = -14'h0006;
         mem[859] =  14'h0031;
         mem[860] = -14'h00e0;
         mem[861] = -14'h003d;
         mem[862] = -14'h0140;
         mem[863] = -14'h0015;
         mem[864] = -14'h007c;
         mem[865] =  14'h002e;
         mem[866] =  14'h009f;
         mem[867] =  14'h00ec;
         mem[868] =  14'h00c6;
         mem[869] = -14'h0116;
         mem[870] = -14'h003b;
         mem[871] =  14'h009e;
         mem[872] =  14'h0102;
         mem[873] =  14'h000b;
         mem[874] =  14'h0001;
         mem[875] =  14'h0004;
         mem[876] = -14'h0049;
         mem[877] = -14'h002a;
         mem[878] = -14'h0002;
         mem[879] = -14'h004b;
         mem[880] = -14'h0007;
         mem[881] = -14'h00b6;
         mem[882] = -14'h0184;
         mem[883] = -14'h0063;
         mem[884] = -14'h0005;
         mem[885] =  14'h0025;
         mem[886] = -14'h0069;
         mem[887] =  14'h0069;
         mem[888] =  14'h008d;
         mem[889] =  14'h0004;
         mem[890] = -14'h004b;
         mem[891] = -14'h0076;
         mem[892] = -14'h0084;
         mem[893] =  14'h0035;
         mem[894] =  14'h016f;
         mem[895] = -14'h000a;
         mem[896] =  14'h0022;
         mem[897] =  14'h001b;
         mem[898] =  14'h0039;
         mem[899] =  14'h0060;
         mem[900] = -14'h0032;
         mem[901] =  14'h0095;
         mem[902] = -14'h00ab;
         mem[903] = -14'h0013;
         mem[904] =  14'h012a;
         mem[905] =  14'h000b;
         mem[906] = -14'h0037;
         mem[907] =  14'h0033;
         mem[908] =  14'h000a;
         mem[909] =  14'h005b;
         mem[910] =  14'h0031;
         mem[911] =  14'h003e;
         mem[912] =  14'h0145;
         mem[913] = -14'h0227;
         mem[914] = -14'h0029;
         mem[915] =  14'h0036;
         mem[916] = -14'h0032;
         mem[917] =  14'h0037;
         mem[918] = -14'h00ff;
         mem[919] =  14'h007d;
         mem[920] = -14'h002c;
         mem[921] = -14'h00bf;
         mem[922] =  14'h008b;
         mem[923] = -14'h0081;
         mem[924] = -14'h00f5;
         mem[925] =  14'h002b;
         mem[926] = -14'h0150;
         mem[927] =  14'h0003;
         mem[928] =  14'h003d;
         mem[929] =  14'h0027;
         mem[930] = -14'h0003;
         mem[931] =  14'h0010;
         mem[932] = -14'h000b;
         mem[933] =  14'h0027;
         mem[934] =  14'h000d;
         mem[935] =  14'h0001;
         mem[936] = -14'h0155;
         mem[937] =  14'h005f;
         mem[938] = -14'h0026;
         mem[939] =  14'h0041;
         mem[940] = -14'h010b;
         mem[941] =  14'h0065;
         mem[942] =  14'h0008;
         mem[943] =  14'h0060;
         mem[944] = -14'h0035;
         mem[945] =  14'h002d;
         mem[946] = -14'h00a5;
         mem[947] = -14'h00fd;
         mem[948] =  14'h0008;
         mem[949] =  14'h0000;
         mem[950] =  14'h0078;
         mem[951] =  14'h0092;
         mem[952] = -14'h01e7;
         mem[953] = -14'h0002;
         mem[954] = -14'h000d;
         mem[955] = -14'h013a;
         mem[956] = -14'h0115;
         mem[957] = -14'h005e;
         mem[958] =  14'h003c;
         mem[959] =  14'h0027;
         mem[960] = -14'h01e6;
         mem[961] =  14'h0005;
         mem[962] =  14'h009c;
         mem[963] =  14'h002f;
         mem[964] =  14'h0226;
         mem[965] =  14'h0021;
         mem[966] = -14'h0084;
         mem[967] =  14'h013c;
         mem[968] = -14'h0008;
         mem[969] =  14'h019b;
         mem[970] = -14'h0001;
         mem[971] =  14'h00f3;
         mem[972] =  14'h01ef;
         mem[973] = -14'h00b2;
         mem[974] =  14'h004e;
         mem[975] =  14'h0092;
         mem[976] =  14'h0094;
         mem[977] =  14'h006e;
         mem[978] = -14'h0033;
         mem[979] =  14'h0119;
         mem[980] =  14'h000e;
         mem[981] = -14'h0055;
         mem[982] =  14'h0039;
         mem[983] =  14'h000f;
         mem[984] =  14'h002f;
         mem[985] = -14'h0042;
         mem[986] =  14'h00b6;
         mem[987] =  14'h0013;
         mem[988] =  14'h00e8;
         mem[989] =  14'h00b9;
         mem[990] =  14'h0035;
         mem[991] = -14'h0003;
         mem[992] = -14'h001d;
         mem[993] = -14'h00c4;
         mem[994] =  14'h000a;
         mem[995] =  14'h0097;
         mem[996] =  14'h0053;
         mem[997] = -14'h0041;
         mem[998] = -14'h008f;
         mem[999] = -14'h0086;
         mem[1000] =  14'h004b;
         mem[1001] =  14'h0040;
         mem[1002] = -14'h0078;
         mem[1003] = -14'h0121;
         mem[1004] = -14'h0043;
         mem[1005] = -14'h0004;
         mem[1006] =  14'h0028;
         mem[1007] = -14'h00b3;
         mem[1008] =  14'h003b;
         mem[1009] =  14'h0074;
         mem[1010] =  14'h0024;
         mem[1011] = -14'h0041;
         mem[1012] = -14'h01c5;
         mem[1013] =  14'h008a;
         mem[1014] =  14'h0055;
         mem[1015] = -14'h012a;
         mem[1016] = -14'h027e;
         mem[1017] =  14'h00f5;
         mem[1018] = -14'h0041;
         mem[1019] = -14'h0102;
         mem[1020] =  14'h0031;
         mem[1021] = -14'h0100;
         mem[1022] =  14'h006a;
         mem[1023] =  14'h0064;
         mem[1024] = -14'h005c;
         mem[1025] =  14'h00ed;
         mem[1026] =  14'h0055;
         mem[1027] =  14'h0017;
         mem[1028] =  14'h003e;
         mem[1029] = -14'h0142;
         mem[1030] =  14'h002b;
         mem[1031] = -14'h00e0;
         mem[1032] =  14'h0021;
         mem[1033] =  14'h0038;
         mem[1034] = -14'h0081;
         mem[1035] =  14'h0075;
         mem[1036] =  14'h008e;
         mem[1037] =  14'h0004;
         mem[1038] = -14'h002b;
         mem[1039] =  14'h0001;
         mem[1040] =  14'h001c;
         mem[1041] = -14'h002f;
         mem[1042] =  14'h00d2;
         mem[1043] = -14'h0058;
         mem[1044] = -14'h0164;
         mem[1045] =  14'h0000;
         mem[1046] =  14'h001d;
         mem[1047] = -14'h0006;
         mem[1048] =  14'h001e;
         mem[1049] = -14'h0035;
         mem[1050] =  14'h0088;
         mem[1051] = -14'h004f;
         mem[1052] = -14'h000d;
         mem[1053] = -14'h0003;
         mem[1054] =  14'h006b;
         mem[1055] =  14'h000a;
         mem[1056] =  14'h00a2;
         mem[1057] =  14'h0002;
         mem[1058] = -14'h0010;
         mem[1059] =  14'h0015;
         mem[1060] = -14'h0066;
         mem[1061] =  14'h0083;
         mem[1062] =  14'h0023;
         mem[1063] =  14'h00a0;
         mem[1064] = -14'h02ba;
         mem[1065] = -14'h0114;
         mem[1066] =  14'h0008;
         mem[1067] =  14'h0070;
         mem[1068] = -14'h003d;
         mem[1069] = -14'h004e;
         mem[1070] =  14'h0042;
         mem[1071] = -14'h01f5;
         mem[1072] =  14'h00bd;
         mem[1073] =  14'h0043;
         mem[1074] =  14'h002b;
         mem[1075] = -14'h0042;
         mem[1076] = -14'h0049;
         mem[1077] = -14'h01c3;
         mem[1078] = -14'h0006;
         mem[1079] =  14'h0107;
         mem[1080] = -14'h013f;
         mem[1081] = -14'h01b7;
         mem[1082] =  14'h0034;
         mem[1083] =  14'h0034;
         mem[1084] =  14'h0033;
         mem[1085] =  14'h01ab;
         mem[1086] = -14'h005a;
         mem[1087] = -14'h002e;
         mem[1088] =  14'h001f;
         mem[1089] = -14'h0128;
         mem[1090] = -14'h04ae;
         mem[1091] = -14'h0025;
         mem[1092] =  14'h0057;
         mem[1093] =  14'h004e;
         mem[1094] =  14'h0006;
         mem[1095] =  14'h0037;
         mem[1096] =  14'h0028;
         mem[1097] = -14'h0002;
         mem[1098] = -14'h00b0;
         mem[1099] =  14'h0137;
         mem[1100] = -14'h0069;
         mem[1101] = -14'h0004;
         mem[1102] =  14'h0031;
         mem[1103] = -14'h006b;
         mem[1104] =  14'h00c8;
         mem[1105] = -14'h0008;
         mem[1106] =  14'h0010;
         mem[1107] = -14'h0030;
         mem[1108] = -14'h00ca;
         mem[1109] =  14'h0096;
         mem[1110] = -14'h004b;
         mem[1111] =  14'h006a;
         mem[1112] =  14'h002b;
         mem[1113] =  14'h0006;
         mem[1114] = -14'h006a;
         mem[1115] =  14'h005b;
         mem[1116] =  14'h00dc;
         mem[1117] =  14'h0019;
         mem[1118] = -14'h00b1;
         mem[1119] =  14'h0009;
         mem[1120] = -14'h00b1;
         mem[1121] = -14'h00f7;
         mem[1122] =  14'h0000;
         mem[1123] = -14'h0053;
         mem[1124] =  14'h00b9;
         mem[1125] =  14'h004d;
         mem[1126] = -14'h001a;
         mem[1127] = -14'h0037;
         mem[1128] = -14'h0028;
         mem[1129] = -14'h0005;
         mem[1130] = -14'h0061;
         mem[1131] = -14'h0045;
         mem[1132] =  14'h0043;
         mem[1133] =  14'h008e;
         mem[1134] =  14'h0007;
         mem[1135] =  14'h0010;
         mem[1136] = -14'h0035;
         mem[1137] =  14'h0010;
         mem[1138] =  14'h0047;
         mem[1139] = -14'h00e2;
         mem[1140] =  14'h0028;
         mem[1141] =  14'h006c;
         mem[1142] =  14'h0028;
         mem[1143] =  14'h001f;
         mem[1144] =  14'h00d2;
         mem[1145] = -14'h002b;
         mem[1146] =  14'h0025;
         mem[1147] = -14'h0007;
         mem[1148] = -14'h00b1;
         mem[1149] = -14'h0006;
         mem[1150] =  14'h0025;
         mem[1151] =  14'h0009;
         mem[1152] =  14'h00cd;
         mem[1153] = -14'h003f;
         mem[1154] =  14'h0032;
         mem[1155] =  14'h0022;
         mem[1156] =  14'h002f;
         mem[1157] = -14'h0059;
         mem[1158] =  14'h0035;
         mem[1159] = -14'h0003;
         mem[1160] = -14'h0074;
         mem[1161] =  14'h0003;
         mem[1162] =  14'h0008;
         mem[1163] =  14'h0045;
         mem[1164] =  14'h002c;
         mem[1165] =  14'h0011;
         mem[1166] =  14'h001e;
         mem[1167] =  14'h011c;
         mem[1168] =  14'h0075;
         mem[1169] = -14'h002f;
         mem[1170] =  14'h0024;
         mem[1171] =  14'h0002;
         mem[1172] = -14'h011a;
         mem[1173] =  14'h0000;
         mem[1174] =  14'h0059;
         mem[1175] = -14'h0007;
         mem[1176] = -14'h0025;
         mem[1177] = -14'h027a;
         mem[1178] = -14'h0070;
         mem[1179] =  14'h00b4;
         mem[1180] =  14'h009d;
         mem[1181] = -14'h0006;
         mem[1182] = -14'h0113;
         mem[1183] = -14'h00b5;
         mem[1184] =  14'h0008;
         mem[1185] =  14'h002c;
         mem[1186] =  14'h0003;
         mem[1187] =  14'h011f;
         mem[1188] =  14'h002c;
         mem[1189] = -14'h002e;
         mem[1190] = -14'h003d;
         mem[1191] =  14'h0000;
         mem[1192] =  14'h0042;
         mem[1193] =  14'h0042;
         mem[1194] =  14'h0096;
         mem[1195] = -14'h0037;
         mem[1196] =  14'h0027;
         mem[1197] = -14'h0122;
         mem[1198] =  14'h013e;
         mem[1199] = -14'h0030;
         mem[1200] =  14'h001f;
         mem[1201] =  14'h0002;
         mem[1202] = -14'h001d;
         mem[1203] = -14'h000e;
         mem[1204] = -14'h000a;
         mem[1205] = -14'h0114;
         mem[1206] =  14'h0000;
         mem[1207] = -14'h00d8;
         mem[1208] = -14'h00cb;
         mem[1209] = -14'h0036;
         mem[1210] =  14'h006d;
         mem[1211] =  14'h0000;
         mem[1212] =  14'h0039;
         mem[1213] = -14'h0062;
         mem[1214] = -14'h00cb;
         mem[1215] =  14'h0068;
         mem[1216] =  14'h00cb;
         mem[1217] =  14'h001d;
         mem[1218] =  14'h0140;
         mem[1219] =  14'h00c5;
         mem[1220] =  14'h0028;
         mem[1221] = -14'h01d7;
         mem[1222] = -14'h0027;
         mem[1223] =  14'h0000;
         mem[1224] =  14'h002b;
         mem[1225] =  14'h0001;
         mem[1226] =  14'h003f;
         mem[1227] = -14'h01d5;
         mem[1228] = -14'h0062;
         mem[1229] =  14'h0005;
         mem[1230] = -14'h0003;
         mem[1231] = -14'h0048;
         mem[1232] = -14'h0168;
         mem[1233] =  14'h00cc;
         mem[1234] = -14'h0015;
         mem[1235] = -14'h0038;
         mem[1236] = -14'h014a;
         mem[1237] =  14'h008b;
         mem[1238] = -14'h0029;
         mem[1239] =  14'h0088;
         mem[1240] = -14'h002b;
         mem[1241] =  14'h000a;
         mem[1242] = -14'h0108;
         mem[1243] =  14'h0051;
         mem[1244] = -14'h01a2;
         mem[1245] = -14'h0033;
         mem[1246] = -14'h00ac;
         mem[1247] =  14'h00e7;
         mem[1248] = -14'h0147;
         mem[1249] =  14'h00c1;
         mem[1250] =  14'h0039;
         mem[1251] =  14'h004f;
         mem[1252] = -14'h0062;
         mem[1253] =  14'h0046;
         mem[1254] = -14'h0136;
         mem[1255] = -14'h004f;
         mem[1256] = -14'h0034;
         mem[1257] =  14'h0034;
         mem[1258] =  14'h0009;
         mem[1259] =  14'h0028;
         mem[1260] =  14'h012e;
         mem[1261] =  14'h0054;
         mem[1262] =  14'h006a;
         mem[1263] =  14'h002d;
         mem[1264] = -14'h0072;
         mem[1265] = -14'h001c;
         mem[1266] = -14'h000a;
         mem[1267] = -14'h000c;
         mem[1268] = -14'h0034;
         mem[1269] = -14'h0122;
         mem[1270] =  14'h0004;
         mem[1271] =  14'h0039;
         mem[1272] =  14'h000a;
         mem[1273] = -14'h011d;
         mem[1274] = -14'h0025;
         mem[1275] = -14'h03f6;
         mem[1276] = -14'h00fc;
         mem[1277] = -14'h00bf;
         mem[1278] =  14'h004d;
         mem[1279] =  14'h0086;
         mem[1280] = -14'h0001;
         mem[1281] =  14'h003c;
         mem[1282] =  14'h0014;
         mem[1283] = -14'h00ab;
         mem[1284] = -14'h0035;
         mem[1285] = -14'h010b;
         mem[1286] =  14'h0000;
         mem[1287] =  14'h009d;
         mem[1288] = -14'h00d9;
         mem[1289] = -14'h0082;
         mem[1290] = -14'h0145;
         mem[1291] =  14'h02b8;
         mem[1292] =  14'h0027;
         mem[1293] =  14'h0023;
         mem[1294] =  14'h0057;
         mem[1295] =  14'h007b;
         mem[1296] = -14'h0202;
         mem[1297] = -14'h001c;
         mem[1298] = -14'h012a;
         mem[1299] =  14'h0024;
         mem[1300] =  14'h009d;
         mem[1301] = -14'h00c0;
         mem[1302] =  14'h0100;
         mem[1303] = -14'h0008;
         mem[1304] = -14'h002f;
         mem[1305] =  14'h004a;
         mem[1306] =  14'h0098;
         mem[1307] =  14'h002d;
         mem[1308] = -14'h0036;
         mem[1309] =  14'h009a;
         mem[1310] = -14'h0006;
         mem[1311] =  14'h0091;
         mem[1312] = -14'h0045;
         mem[1313] =  14'h003f;
         mem[1314] = -14'h0034;
         mem[1315] = -14'h00c2;
         mem[1316] = -14'h0041;
         mem[1317] = -14'h0049;
         mem[1318] =  14'h0008;
         mem[1319] = -14'h0044;
         mem[1320] = -14'h0125;
         mem[1321] =  14'h004c;
         mem[1322] = -14'h0153;
         mem[1323] =  14'h00b4;
         mem[1324] = -14'h0073;
         mem[1325] = -14'h000f;
         mem[1326] =  14'h0070;
         mem[1327] =  14'h00b4;
         mem[1328] =  14'h003d;
         mem[1329] =  14'h001d;
         mem[1330] = -14'h0118;
         mem[1331] =  14'h0013;
         mem[1332] =  14'h001d;
         mem[1333] =  14'h002a;
         mem[1334] = -14'h00da;
         mem[1335] =  14'h006b;
         mem[1336] = -14'h00a6;
         mem[1337] =  14'h0027;
         mem[1338] = -14'h0057;
         mem[1339] =  14'h00ca;
         mem[1340] = -14'h0039;
         mem[1341] = -14'h0001;
         mem[1342] = -14'h000f;
         mem[1343] =  14'h0033;
         mem[1344] = -14'h0039;
         mem[1345] =  14'h003f;
         mem[1346] =  14'h00ba;
         mem[1347] =  14'h0049;
         mem[1348] = -14'h011d;
         mem[1349] =  14'h00aa;
         mem[1350] = -14'h0043;
         mem[1351] =  14'h0030;
         mem[1352] = -14'h0119;
         mem[1353] = -14'h02ee;
         mem[1354] = -14'h0046;
         mem[1355] = -14'h00a0;
         mem[1356] = -14'h005e;
         mem[1357] =  14'h0031;
         mem[1358] = -14'h01f2;
         mem[1359] =  14'h002f;
         mem[1360] = -14'h0027;
         mem[1361] =  14'h001c;
         mem[1362] =  14'h0005;
         mem[1363] =  14'h00fc;
         mem[1364] = -14'h000b;
         mem[1365] = -14'h012d;
         mem[1366] = -14'h00ef;
         mem[1367] = -14'h017f;
         mem[1368] =  14'h0190;
         mem[1369] = -14'h00ad;
         mem[1370] =  14'h001b;
         mem[1371] =  14'h0007;
         mem[1372] = -14'h002b;
         mem[1373] =  14'h0021;
         mem[1374] = -14'h0085;
         mem[1375] =  14'h0021;
         mem[1376] =  14'h007c;
         mem[1377] =  14'h0002;
         mem[1378] =  14'h008a;
         mem[1379] = -14'h0005;
         mem[1380] =  14'h007f;
         mem[1381] = -14'h0038;
         mem[1382] =  14'h0004;
         mem[1383] =  14'h0012;
         mem[1384] = -14'h0002;
         mem[1385] = -14'h0049;
         mem[1386] = -14'h023b;
         mem[1387] =  14'h0068;
         mem[1388] = -14'h0033;
         mem[1389] =  14'h0045;
         mem[1390] =  14'h0016;
         mem[1391] = -14'h0118;
         mem[1392] = -14'h0025;
         mem[1393] = -14'h006c;
         mem[1394] = -14'h0034;
         mem[1395] =  14'h0007;
         mem[1396] = -14'h0037;
         mem[1397] =  14'h0024;
         mem[1398] = -14'h0003;
         mem[1399] =  14'h0020;
         mem[1400] = -14'h00a2;
         mem[1401] = -14'h0078;
         mem[1402] =  14'h01f3;
         mem[1403] = -14'h021e;
         mem[1404] =  14'h007e;
         mem[1405] =  14'h00c3;
         mem[1406] =  14'h0065;
         mem[1407] = -14'h00a2;
         mem[1408] = -14'h0093;
         mem[1409] = -14'h00af;
         mem[1410] =  14'h0046;
         mem[1411] =  14'h003e;
         mem[1412] =  14'h0045;
         mem[1413] =  14'h001d;
         mem[1414] =  14'h003d;
         mem[1415] = -14'h00a9;
         mem[1416] =  14'h006b;
         mem[1417] = -14'h0030;
         mem[1418] = -14'h00ea;
         mem[1419] =  14'h0064;
         mem[1420] =  14'h0071;
         mem[1421] =  14'h0000;
         mem[1422] =  14'h002b;
         mem[1423] = -14'h00cd;
         mem[1424] =  14'h002e;
         mem[1425] = -14'h0035;
         mem[1426] =  14'h0038;
         mem[1427] = -14'h0030;
         mem[1428] =  14'h0025;
         mem[1429] = -14'h003c;
         mem[1430] =  14'h0037;
         mem[1431] = -14'h009a;
         mem[1432] =  14'h0027;
         mem[1433] =  14'h0003;
         mem[1434] = -14'h0017;
         mem[1435] = -14'h0166;
         mem[1436] = -14'h007e;
         mem[1437] = -14'h0003;
         mem[1438] =  14'h0000;
         mem[1439] = -14'h004b;
         mem[1440] =  14'h0033;
         mem[1441] =  14'h000c;
         mem[1442] =  14'h0026;
         mem[1443] = -14'h0043;
         mem[1444] =  14'h010a;
         mem[1445] = -14'h012d;
         mem[1446] = -14'h000e;
         mem[1447] = -14'h003e;
         mem[1448] =  14'h002b;
         mem[1449] = -14'h0111;
         mem[1450] = -14'h0156;
         mem[1451] =  14'h0074;
         mem[1452] = -14'h005f;
         mem[1453] =  14'h0004;
         mem[1454] =  14'h003c;
         mem[1455] = -14'h0052;
         mem[1456] = -14'h0105;
         mem[1457] = -14'h002c;
         mem[1458] =  14'h003d;
         mem[1459] = -14'h0035;
         mem[1460] =  14'h002c;
         mem[1461] = -14'h0008;
         mem[1462] =  14'h0101;
         mem[1463] = -14'h0099;
         mem[1464] =  14'h0060;
         mem[1465] = -14'h00b7;
         mem[1466] =  14'h0052;
         mem[1467] = -14'h00c6;
         mem[1468] = -14'h000f;
         mem[1469] =  14'h0093;
         mem[1470] =  14'h0020;
         mem[1471] = -14'h000d;
         mem[1472] = -14'h00a2;
         mem[1473] = -14'h002e;
         mem[1474] = -14'h021f;
         mem[1475] =  14'h0016;
         mem[1476] =  14'h0004;
         mem[1477] = -14'h011a;
         mem[1478] = -14'h0062;
         mem[1479] = -14'h002b;
         mem[1480] = -14'h0062;
         mem[1481] =  14'h005a;
         mem[1482] = -14'h00e9;
         mem[1483] = -14'h0005;
         mem[1484] =  14'h0000;
         mem[1485] =  14'h0058;
         mem[1486] =  14'h0059;
         mem[1487] =  14'h000a;
         mem[1488] = -14'h000d;
         mem[1489] = -14'h0052;
         mem[1490] =  14'h0a00;
         mem[1491] =  14'h0055;
         mem[1492] =  14'h002d;
         mem[1493] =  14'h002a;
         mem[1494] = -14'h018a;
         mem[1495] = -14'h00ff;
         mem[1496] =  14'h0003;
         mem[1497] = -14'h0033;
         mem[1498] =  14'h0115;
         mem[1499] =  14'h0032;
         mem[1500] =  14'h0011;
         mem[1501] = -14'h00d7;
         mem[1502] =  14'h005d;
         mem[1503] = -14'h0046;
         mem[1504] =  14'h001b;
         mem[1505] = -14'h003b;
         mem[1506] =  14'h002c;
         mem[1507] = -14'h00d6;
         mem[1508] = -14'h002c;
         mem[1509] = -14'h0025;
         mem[1510] =  14'h0003;
         mem[1511] = -14'h00c2;
         mem[1512] =  14'h00c3;
         mem[1513] = -14'h0002;
         mem[1514] =  14'h0038;
         mem[1515] = -14'h005b;
         mem[1516] =  14'h0042;
         mem[1517] =  14'h0007;
         mem[1518] = -14'h00ab;
         mem[1519] = -14'h0025;
         mem[1520] =  14'h0035;
         mem[1521] =  14'h000c;
         mem[1522] =  14'h0021;
         mem[1523] =  14'h0066;
         mem[1524] = -14'h00b6;
         mem[1525] = -14'h004a;
         mem[1526] =  14'h0000;
         mem[1527] = -14'h0002;
         mem[1528] = -14'h012d;
         mem[1529] = -14'h01db;
         mem[1530] =  14'h0063;
         mem[1531] = -14'h011c;
         mem[1532] =  14'h00fc;
         mem[1533] = -14'h00b1;
         mem[1534] =  14'h0011;
         mem[1535] = -14'h027f;
         mem[1536] =  14'h0026;
         mem[1537] = -14'h0223;
         mem[1538] =  14'h00c8;
         mem[1539] = -14'h00b8;
         mem[1540] = -14'h015d;
         mem[1541] =  14'h00ba;
         mem[1542] =  14'h0031;
         mem[1543] = -14'h000a;
         mem[1544] =  14'h0000;
         mem[1545] = -14'h01d1;
         mem[1546] =  14'h0035;
         mem[1547] = -14'h016a;
         mem[1548] = -14'h001e;
         mem[1549] =  14'h0042;
         mem[1550] =  14'h002c;
         mem[1551] = -14'h009c;
         mem[1552] =  14'h004d;
         mem[1553] = -14'h003a;
         mem[1554] =  14'h0035;
         mem[1555] =  14'h0011;
         mem[1556] =  14'h0085;
         mem[1557] = -14'h007e;
         mem[1558] =  14'h0014;
         mem[1559] =  14'h0080;
         mem[1560] = -14'h0095;
         mem[1561] =  14'h0099;
         mem[1562] =  14'h0037;
         mem[1563] =  14'h009c;
         mem[1564] =  14'h0081;
         mem[1565] =  14'h0069;
         mem[1566] =  14'h0018;
         mem[1567] =  14'h003c;
         mem[1568] =  14'h002e;
         mem[1569] =  14'h000a;
         mem[1570] = -14'h00d1;
         mem[1571] =  14'h0039;
         mem[1572] = -14'h0032;
         mem[1573] =  14'h00ce;
         mem[1574] =  14'h0005;
         mem[1575] = -14'h0013;
         mem[1576] =  14'h006c;
         mem[1577] =  14'h0027;
         mem[1578] =  14'h0002;
         mem[1579] = -14'h00e8;
         mem[1580] = -14'h0042;
         mem[1581] =  14'h0044;
         mem[1582] =  14'h0019;
         mem[1583] =  14'h0039;
         mem[1584] = -14'h0043;
         mem[1585] =  14'h0023;
         mem[1586] = -14'h00b9;
         mem[1587] =  14'h0083;
         mem[1588] = -14'h0115;
         mem[1589] =  14'h0025;
         mem[1590] =  14'h0007;
         mem[1591] =  14'h0040;
         mem[1592] =  14'h0077;
         mem[1593] =  14'h0021;
         mem[1594] = -14'h003d;
         mem[1595] = -14'h009d;
         mem[1596] =  14'h0008;
         mem[1597] =  14'h002c;
         mem[1598] = -14'h0046;
         mem[1599] =  14'h003d;
         mem[1600] =  14'h0024;
         mem[1601] = -14'h003d;
         mem[1602] = -14'h00f2;
         mem[1603] =  14'h0018;
         mem[1604] = -14'h00dc;
         mem[1605] =  14'h0062;
         mem[1606] =  14'h0007;
         mem[1607] =  14'h000c;
         mem[1608] = -14'h003d;
         mem[1609] =  14'h0040;
         mem[1610] = -14'h003b;
         mem[1611] = -14'h0034;
         mem[1612] = -14'h000a;
         mem[1613] =  14'h009a;
         mem[1614] =  14'h00e5;
         mem[1615] = -14'h0045;
         mem[1616] =  14'h0005;
         mem[1617] =  14'h00a3;
         mem[1618] = -14'h003b;
         mem[1619] =  14'h0008;
         mem[1620] =  14'h0008;
         mem[1621] =  14'h002a;
         mem[1622] = -14'h01fc;
         mem[1623] =  14'h0061;
         mem[1624] = -14'h00eb;
         mem[1625] =  14'h003a;
         mem[1626] =  14'h008a;
         mem[1627] = -14'h0020;
         mem[1628] =  14'h0052;
         mem[1629] = -14'h009b;
         mem[1630] = -14'h0007;
         mem[1631] =  14'h0007;
         mem[1632] = -14'h000b;
         mem[1633] =  14'h0002;
         mem[1634] = -14'h0026;
         mem[1635] =  14'h002b;
         mem[1636] =  14'h0079;
         mem[1637] = -14'h0059;
         mem[1638] = -14'h000a;
         mem[1639] =  14'h0028;
         mem[1640] = -14'h0033;
         mem[1641] =  14'h0016;
         mem[1642] = -14'h0001;
         mem[1643] =  14'h0024;
         mem[1644] =  14'h0001;
         mem[1645] =  14'h0026;
         mem[1646] = -14'h0073;
         mem[1647] =  14'h0047;
         mem[1648] =  14'h00ac;
         mem[1649] =  14'h0017;
         mem[1650] =  14'h0055;
         mem[1651] =  14'h0023;
         mem[1652] = -14'h00ae;
         mem[1653] =  14'h008a;
         mem[1654] =  14'h00c9;
         mem[1655] = -14'h007a;
         mem[1656] = -14'h009c;
         mem[1657] =  14'h006a;
         mem[1658] =  14'h00bd;
         mem[1659] = -14'h0022;
         mem[1660] =  14'h009d;
         mem[1661] =  14'h0025;
         mem[1662] = -14'h0117;
         mem[1663] =  14'h0039;
         mem[1664] =  14'h000e;
         mem[1665] = -14'h0036;
         mem[1666] =  14'h009e;
         mem[1667] =  14'h0040;
         mem[1668] =  14'h000a;
         mem[1669] =  14'h0000;
         mem[1670] = -14'h0056;
         mem[1671] =  14'h0002;
         mem[1672] =  14'h007b;
         mem[1673] = -14'h002c;
         mem[1674] =  14'h0002;
         mem[1675] =  14'h0051;
         mem[1676] = -14'h002c;
         mem[1677] = -14'h0002;
         mem[1678] =  14'h0079;
         mem[1679] = -14'h0044;
         mem[1680] = -14'h0105;
         mem[1681] =  14'h0092;
         mem[1682] = -14'h006b;
         mem[1683] =  14'h02e1;
         mem[1684] =  14'h0216;
         mem[1685] =  14'h0024;
         mem[1686] =  14'h008a;
         mem[1687] = -14'h0190;
         mem[1688] = -14'h0025;
         mem[1689] =  14'h0021;
         mem[1690] = -14'h000e;
         mem[1691] =  14'h0093;
         mem[1692] =  14'h0005;
         mem[1693] =  14'h005f;
         mem[1694] = -14'h003a;
         mem[1695] = -14'h0068;
         mem[1696] = -14'h01b1;
         mem[1697] = -14'h0075;
         mem[1698] =  14'h0027;
         mem[1699] =  14'h0008;
         mem[1700] = -14'h002f;
         mem[1701] = -14'h007a;
         mem[1702] = -14'h0043;
         mem[1703] =  14'h000d;
         mem[1704] = -14'h0022;
         mem[1705] = -14'h00ad;
         mem[1706] = -14'h00bb;
         mem[1707] =  14'h004e;
         mem[1708] = -14'h0008;
         mem[1709] =  14'h0053;
         mem[1710] =  14'h006f;
         mem[1711] = -14'h04c2;
         mem[1712] = -14'h000f;
         mem[1713] = -14'h0008;
         mem[1714] = -14'h00c4;
         mem[1715] = -14'h0015;
         mem[1716] = -14'h0006;
         mem[1717] = -14'h023a;
         mem[1718] = -14'h003d;
         mem[1719] =  14'h0020;
         mem[1720] = -14'h0032;
         mem[1721] =  14'h0023;
         mem[1722] =  14'h0007;
         mem[1723] = -14'h0024;
         mem[1724] = -14'h000c;
         mem[1725] = -14'h0011;
         mem[1726] = -14'h000a;
         mem[1727] =  14'h00d1;
         mem[1728] = -14'h0030;
         mem[1729] =  14'h009b;
         mem[1730] =  14'h0070;
         mem[1731] =  14'h008c;
         mem[1732] =  14'h0076;
         mem[1733] = -14'h00fb;
         mem[1734] =  14'h00b6;
         mem[1735] = -14'h0037;
         mem[1736] =  14'h0040;
         mem[1737] = -14'h0114;
         mem[1738] =  14'h0083;
         mem[1739] = -14'h013e;
         mem[1740] =  14'h0034;
         mem[1741] = -14'h0059;
         mem[1742] =  14'h0034;
         mem[1743] =  14'h0005;
         mem[1744] =  14'h008c;
         mem[1745] =  14'h0044;
         mem[1746] = -14'h0105;
         mem[1747] = -14'h00df;
         mem[1748] =  14'h00cd;
         mem[1749] =  14'h003a;
         mem[1750] =  14'h0024;
         mem[1751] = -14'h01e9;
         mem[1752] = -14'h0053;
         mem[1753] =  14'h0000;
         mem[1754] =  14'h002a;
         mem[1755] =  14'h00d5;
         mem[1756] = -14'h0012;
         mem[1757] = -14'h0127;
         mem[1758] =  14'h0026;
         mem[1759] =  14'h0081;
         mem[1760] =  14'h004a;
         mem[1761] = -14'h00e4;
         mem[1762] = -14'h000b;
         mem[1763] = -14'h0005;
         mem[1764] =  14'h00f7;
         mem[1765] = -14'h002c;
         mem[1766] =  14'h0046;
         mem[1767] = -14'h01c7;
         mem[1768] = -14'h0006;
         mem[1769] = -14'h00b4;
         mem[1770] =  14'h0054;
         mem[1771] = -14'h004d;
         mem[1772] =  14'h0094;
         mem[1773] =  14'h000b;
         mem[1774] =  14'h0030;
         mem[1775] = -14'h00b0;
         mem[1776] =  14'h0027;
         mem[1777] = -14'h0099;
         mem[1778] =  14'h0060;
         mem[1779] =  14'h0084;
         mem[1780] =  14'h0024;
         mem[1781] =  14'h012e;
         mem[1782] =  14'h00ea;
         mem[1783] = -14'h000e;
         mem[1784] = -14'h0100;
         mem[1785] = -14'h0001;
         mem[1786] = -14'h01af;
         mem[1787] = -14'h0027;
         mem[1788] = -14'h002f;
         mem[1789] = -14'h0004;
         mem[1790] = -14'h0041;
         mem[1791] = -14'h004f;
         mem[1792] =  14'h006b;
         mem[1793] =  14'h00ed;
         mem[1794] =  14'h0067;
         mem[1795] = -14'h00fd;
         mem[1796] =  14'h0041;
         mem[1797] =  14'h001e;
         mem[1798] = -14'h0107;
         mem[1799] =  14'h0008;
         mem[1800] =  14'h0000;
         mem[1801] = -14'h0057;
         mem[1802] =  14'h0026;
         mem[1803] =  14'h0007;
         mem[1804] =  14'h002f;
         mem[1805] =  14'h0014;
         mem[1806] =  14'h0039;
         mem[1807] =  14'h0010;
         mem[1808] =  14'h0038;
         mem[1809] = -14'h006f;
         mem[1810] =  14'h0061;
         mem[1811] =  14'h0066;
         mem[1812] = -14'h0044;
         mem[1813] = -14'h0011;
         mem[1814] =  14'h0028;
         mem[1815] =  14'h00c6;
         mem[1816] = -14'h009a;
         mem[1817] = -14'h009e;
         mem[1818] = -14'h00b5;
         mem[1819] = -14'h0012;
         mem[1820] =  14'h0015;
         mem[1821] =  14'h0046;
         mem[1822] = -14'h000f;
         mem[1823] = -14'h000f;
         mem[1824] =  14'h0081;
         mem[1825] =  14'h004e;
         mem[1826] = -14'h0080;
         mem[1827] =  14'h0064;
         mem[1828] =  14'h0033;
         mem[1829] = -14'h0088;
         mem[1830] = -14'h00a0;
         mem[1831] =  14'h016b;
         mem[1832] =  14'h0028;
         mem[1833] = -14'h002a;
         mem[1834] =  14'h0026;
         mem[1835] =  14'h006c;
         mem[1836] =  14'h0025;
         mem[1837] =  14'h0044;
         mem[1838] =  14'h006e;
         mem[1839] =  14'h00b1;
         mem[1840] = -14'h0056;
         mem[1841] = -14'h015a;
         mem[1842] = -14'h000f;
         mem[1843] = -14'h000a;
         mem[1844] =  14'h003c;
         mem[1845] = -14'h0036;
         mem[1846] =  14'h0035;
         mem[1847] = -14'h0002;
         mem[1848] =  14'h000b;
         mem[1849] = -14'h003c;
         mem[1850] =  14'h0046;
         mem[1851] =  14'h0013;
         mem[1852] = -14'h0005;
         mem[1853] = -14'h000a;
         mem[1854] =  14'h0080;
         mem[1855] =  14'h0043;
         mem[1856] =  14'h0051;
         mem[1857] = -14'h0023;
         mem[1858] = -14'h0007;
         mem[1859] = -14'h0003;
         mem[1860] =  14'h000b;
         mem[1861] =  14'h0051;
         mem[1862] =  14'h002b;
         mem[1863] = -14'h0025;
         mem[1864] =  14'h001f;
         mem[1865] = -14'h0006;
         mem[1866] =  14'h002a;
         mem[1867] =  14'h0120;
         mem[1868] =  14'h0009;
         mem[1869] = -14'h0034;
         mem[1870] =  14'h008a;
         mem[1871] =  14'h0000;
         mem[1872] =  14'h006b;
         mem[1873] =  14'h0020;
         mem[1874] =  14'h0037;
         mem[1875] = -14'h0069;
         mem[1876] =  14'h001c;
         mem[1877] = -14'h004c;
         mem[1878] =  14'h003f;
         mem[1879] = -14'h003b;
         mem[1880] =  14'h0027;
         mem[1881] = -14'h000d;
         mem[1882] = -14'h0253;
         mem[1883] = -14'h0002;
         mem[1884] = -14'h00ab;
         mem[1885] = -14'h0144;
         mem[1886] =  14'h0003;
         mem[1887] = -14'h0006;
         mem[1888] = -14'h0007;
         mem[1889] = -14'h0024;
         mem[1890] =  14'h0060;
         mem[1891] = -14'h0363;
         mem[1892] =  14'h0004;
         mem[1893] = -14'h002d;
         mem[1894] = -14'h004f;
         mem[1895] =  14'h0054;
         mem[1896] = -14'h002e;
         mem[1897] = -14'h0121;
         mem[1898] =  14'h0011;
         mem[1899] = -14'h0004;
         mem[1900] = -14'h002f;
         mem[1901] = -14'h0004;
         mem[1902] =  14'h0003;
         mem[1903] = -14'h006a;
         mem[1904] =  14'h001e;
         mem[1905] = -14'h0032;
         mem[1906] = -14'h0006;
         mem[1907] = -14'h0006;
         mem[1908] =  14'h0010;
         mem[1909] =  14'h0000;
         mem[1910] =  14'h007d;
         mem[1911] =  14'h0082;
         mem[1912] = -14'h0029;
         mem[1913] = -14'h0121;
         mem[1914] =  14'h0016;
         mem[1915] = -14'h0025;
         mem[1916] =  14'h00db;
         mem[1917] =  14'h0056;
         mem[1918] =  14'h001e;
         mem[1919] = -14'h003e;
         mem[1920] = -14'h004b;
         mem[1921] =  14'h0000;
         mem[1922] = -14'h0024;
         mem[1923] = -14'h0048;
         mem[1924] = -14'h0048;
         mem[1925] =  14'h009c;
         mem[1926] = -14'h0069;
         mem[1927] =  14'h004b;
         mem[1928] =  14'h0024;
         mem[1929] = -14'h00af;
         mem[1930] =  14'h001f;
         mem[1931] = -14'h0106;
         mem[1932] =  14'h0036;
         mem[1933] =  14'h007c;
         mem[1934] =  14'h0050;
         mem[1935] = -14'h004c;
         mem[1936] = -14'h00ff;
         mem[1937] =  14'h0005;
         mem[1938] = -14'h0007;
         mem[1939] = -14'h0044;
         mem[1940] = -14'h0060;
         mem[1941] =  14'h0069;
         mem[1942] =  14'h0021;
         mem[1943] =  14'h0000;
         mem[1944] = -14'h0036;
         mem[1945] = -14'h0002;
         mem[1946] = -14'h000e;
         mem[1947] = -14'h00bb;
         mem[1948] =  14'h002a;
         mem[1949] = -14'h00ee;
         mem[1950] =  14'h0040;
         mem[1951] =  14'h0011;
         mem[1952] =  14'h0029;
         mem[1953] = -14'h0005;
         mem[1954] = -14'h0027;
         mem[1955] =  14'h00bc;
         mem[1956] =  14'h002e;
         mem[1957] = -14'h0003;
         mem[1958] = -14'h0009;
         mem[1959] =  14'h006c;
         mem[1960] = -14'h00fc;
         mem[1961] =  14'h0036;
         mem[1962] =  14'h004c;
         mem[1963] = -14'h003e;
         mem[1964] =  14'h0024;
         mem[1965] = -14'h0034;
         mem[1966] =  14'h0066;
         mem[1967] = -14'h000d;
         mem[1968] =  14'h013e;
         mem[1969] =  14'h0099;
         mem[1970] =  14'h0028;
         mem[1971] = -14'h0074;
         mem[1972] =  14'h0039;
         mem[1973] = -14'h003d;
         mem[1974] =  14'h000a;
         mem[1975] =  14'h0024;
         mem[1976] =  14'h0015;
         mem[1977] = -14'h0008;
         mem[1978] =  14'h000d;
         mem[1979] = -14'h0056;
         mem[1980] = -14'h0068;
         mem[1981] = -14'h00d1;
         mem[1982] = -14'h0053;
         mem[1983] =  14'h000b;
         mem[1984] =  14'h0038;
         mem[1985] = -14'h0038;
         mem[1986] =  14'h002d;
         mem[1987] = -14'h00df;
         mem[1988] =  14'h0005;
         mem[1989] =  14'h000d;
         mem[1990] =  14'h0058;
         mem[1991] = -14'h00a7;
         mem[1992] =  14'h0096;
         mem[1993] = -14'h0052;
         mem[1994] = -14'h003c;
         mem[1995] = -14'h019b;
         mem[1996] =  14'h0026;
         mem[1997] =  14'h0003;
         mem[1998] =  14'h008e;
         mem[1999] = -14'h0060;
         mem[2000] = -14'h006d;
         mem[2001] =  14'h000b;
         mem[2002] =  14'h000b;
         mem[2003] = -14'h002d;
         mem[2004] = -14'h004c;
         mem[2005] = -14'h000c;
         mem[2006] =  14'h002f;
         mem[2007] = -14'h002e;
         mem[2008] = -14'h0010;
         mem[2009] = -14'h000f;
         mem[2010] = -14'h0169;
         mem[2011] = -14'h000d;
         mem[2012] =  14'h0071;
         mem[2013] = -14'h002f;
         mem[2014] =  14'h00d0;
         mem[2015] =  14'h0000;
         mem[2016] =  14'h000e;
         mem[2017] = -14'h0033;
         mem[2018] =  14'h003a;
         mem[2019] = -14'h0042;
         mem[2020] =  14'h0021;
         mem[2021] =  14'h0004;
         mem[2022] =  14'h0024;
         mem[2023] = -14'h008f;
         mem[2024] = -14'h004b;
         mem[2025] =  14'h0003;
         mem[2026] =  14'h0000;
         mem[2027] = -14'h000a;
         mem[2028] = -14'h0040;
         mem[2029] = -14'h002e;
         mem[2030] =  14'h0025;
         mem[2031] =  14'h0057;
         mem[2032] = -14'h0102;
         mem[2033] =  14'h0015;
         mem[2034] =  14'h000f;
         mem[2035] =  14'h0015;
         mem[2036] =  14'h001e;
         mem[2037] =  14'h01e6;
         mem[2038] =  14'h0042;
         mem[2039] =  14'h000b;
         mem[2040] = -14'h000a;
         mem[2041] = -14'h0012;
         mem[2042] =  14'h00dc;
         mem[2043] = -14'h0028;
         mem[2044] = -14'h028e;
         mem[2045] = -14'h00b5;
         mem[2046] =  14'h01a6;
         mem[2047] = -14'h002c;
         mem[2048] = -14'h0014;
         mem[2049] =  14'h0019;
         mem[2050] =  14'h0044;
         mem[2051] = -14'h00d9;
         mem[2052] = -14'h008f;
         mem[2053] =  14'h00f8;
         mem[2054] = -14'h0119;
         mem[2055] =  14'h00d2;
         mem[2056] =  14'h0049;
         mem[2057] = -14'h00c8;
         mem[2058] =  14'h0034;
         mem[2059] =  14'h0010;
         mem[2060] = -14'h002d;
         mem[2061] =  14'h011b;
         mem[2062] =  14'h00b2;
         mem[2063] = -14'h0040;
         mem[2064] =  14'h001d;
         mem[2065] = -14'h000d;
         mem[2066] =  14'h000b;
         mem[2067] = -14'h0058;
         mem[2068] =  14'h001d;
         mem[2069] = -14'h0070;
         mem[2070] = -14'h00ba;
         mem[2071] = -14'h002e;
         mem[2072] =  14'h0009;
         mem[2073] = -14'h0035;
         mem[2074] =  14'h0047;
         mem[2075] =  14'h008b;
         mem[2076] = -14'h001c;
         mem[2077] = -14'h002a;
         mem[2078] = -14'h00c9;
         mem[2079] =  14'h00aa;
         mem[2080] =  14'h0029;
         mem[2081] = -14'h0028;
         mem[2082] = -14'h047d;
         mem[2083] =  14'h0003;
         mem[2084] =  14'h0021;
         mem[2085] = -14'h00bb;
         mem[2086] =  14'h0023;
         mem[2087] =  14'h0014;
         mem[2088] =  14'h006b;
         mem[2089] =  14'h00a5;
         mem[2090] =  14'h0024;
         mem[2091] = -14'h0257;
         mem[2092] =  14'h0015;
         mem[2093] = -14'h000d;
         mem[2094] =  14'h00bc;
         mem[2095] =  14'h00b2;
         mem[2096] = -14'h0034;
         mem[2097] = -14'h002d;
         mem[2098] =  14'h0030;
         mem[2099] =  14'h0347;
         mem[2100] =  14'h003c;
         mem[2101] =  14'h004c;
         mem[2102] = -14'h0022;
         mem[2103] = -14'h004a;
         mem[2104] = -14'h00ae;
         mem[2105] = -14'h0003;
         mem[2106] =  14'h0116;
         mem[2107] =  14'h0032;
         mem[2108] = -14'h0091;
         mem[2109] =  14'h0024;
         mem[2110] = -14'h008e;
         mem[2111] = -14'h003a;
         mem[2112] =  14'h0032;
         mem[2113] = -14'h0057;
         mem[2114] =  14'h0017;
         mem[2115] =  14'h0000;
         mem[2116] =  14'h0006;
         mem[2117] = -14'h000c;
         mem[2118] = -14'h0083;
         mem[2119] = -14'h0131;
         mem[2120] =  14'h0009;
         mem[2121] =  14'h007e;
         mem[2122] =  14'h0066;
         mem[2123] =  14'h00b0;
         mem[2124] =  14'h0041;
         mem[2125] =  14'h004f;
         mem[2126] = -14'h0046;
         mem[2127] = -14'h0045;
         mem[2128] = -14'h00e2;
         mem[2129] = -14'h008b;
         mem[2130] =  14'h0006;
         mem[2131] =  14'h0036;
         mem[2132] = -14'h00ae;
         mem[2133] =  14'h003c;
         mem[2134] = -14'h0036;
         mem[2135] =  14'h00ac;
         mem[2136] = -14'h00ce;
         mem[2137] =  14'h0004;
         mem[2138] =  14'h0078;
         mem[2139] = -14'h000f;
         mem[2140] = -14'h0104;
         mem[2141] =  14'h0001;
         mem[2142] =  14'h0000;
         mem[2143] =  14'h003f;
         mem[2144] = -14'h00f0;
         mem[2145] =  14'h0002;
         mem[2146] = -14'h005b;
         mem[2147] = -14'h01a1;
         mem[2148] = -14'h01b2;
         mem[2149] =  14'h0084;
         mem[2150] =  14'h00f3;
         mem[2151] = -14'h0128;
         mem[2152] = -14'h0054;
         mem[2153] =  14'h0000;
         mem[2154] = -14'h00c6;
         mem[2155] =  14'h00be;
         mem[2156] = -14'h002f;
         mem[2157] =  14'h0008;
         mem[2158] = -14'h0147;
         mem[2159] =  14'h00aa;
         mem[2160] = -14'h0005;
         mem[2161] =  14'h003b;
         mem[2162] =  14'h00db;
         mem[2163] =  14'h0007;
         mem[2164] = -14'h00f7;
         mem[2165] =  14'h0084;
         mem[2166] = -14'h002e;
         mem[2167] =  14'h0051;
         mem[2168] = -14'h000f;
         mem[2169] =  14'h0005;
         mem[2170] = -14'h004a;
         mem[2171] =  14'h003b;
         mem[2172] = -14'h0042;
         mem[2173] =  14'h000f;
         mem[2174] =  14'h01a3;
         mem[2175] = -14'h0072;
         mem[2176] = -14'h003c;
         mem[2177] =  14'h00ce;
         mem[2178] = -14'h0054;
         mem[2179] = -14'h016b;
         mem[2180] =  14'h0095;
         mem[2181] =  14'h0063;
         mem[2182] = -14'h0028;
         mem[2183] =  14'h0002;
         mem[2184] = -14'h0008;
         mem[2185] =  14'h0029;
         mem[2186] =  14'h008b;
         mem[2187] = -14'h0003;
         mem[2188] =  14'h00c2;
         mem[2189] = -14'h00bd;
         mem[2190] =  14'h0189;
         mem[2191] =  14'h0034;
         mem[2192] =  14'h000d;
         mem[2193] =  14'h004b;
         mem[2194] = -14'h0048;
         mem[2195] =  14'h0016;
         mem[2196] =  14'h0040;
         mem[2197] =  14'h0004;
         mem[2198] = -14'h0040;
         mem[2199] =  14'h0016;
         mem[2200] = -14'h0068;
         mem[2201] =  14'h002c;
         mem[2202] = -14'h0009;
         mem[2203] = -14'h00ce;
         mem[2204] = -14'h002c;
         mem[2205] = -14'h01f7;
         mem[2206] = -14'h0107;
         mem[2207] =  14'h001f;
         mem[2208] =  14'h00be;
         mem[2209] = -14'h0071;
         mem[2210] = -14'h002c;
         mem[2211] = -14'h001f;
         mem[2212] = -14'h0055;
         mem[2213] =  14'h0025;
         mem[2214] = -14'h0007;
         mem[2215] =  14'h0054;
         mem[2216] = -14'h00d5;
         mem[2217] =  14'h002d;
         mem[2218] =  14'h0011;
         mem[2219] = -14'h0060;
         mem[2220] = -14'h0035;
         mem[2221] =  14'h0074;
         mem[2222] =  14'h0013;
         mem[2223] = -14'h0048;
         mem[2224] = -14'h008d;
         mem[2225] = -14'h0035;
         mem[2226] =  14'h0011;
         mem[2227] =  14'h00c1;
         mem[2228] = -14'h0051;
         mem[2229] = -14'h0123;
         mem[2230] =  14'h0030;
         mem[2231] =  14'h002a;
         mem[2232] = -14'h0005;
         mem[2233] =  14'h0087;
         mem[2234] = -14'h0047;
         mem[2235] =  14'h0010;
         mem[2236] =  14'h0082;
         mem[2237] = -14'h0173;
         mem[2238] =  14'h0006;
         mem[2239] =  14'h001e;
         mem[2240] = -14'h0105;
         mem[2241] =  14'h002f;
         mem[2242] = -14'h00d4;
         mem[2243] =  14'h0024;
         mem[2244] =  14'h007a;
         mem[2245] = -14'h009c;
         mem[2246] =  14'h001e;
         mem[2247] =  14'h0010;
         mem[2248] = -14'h0024;
         mem[2249] =  14'h0010;
         mem[2250] = -14'h008a;
         mem[2251] =  14'h0064;
         mem[2252] = -14'h008a;
         mem[2253] =  14'h0009;
         mem[2254] =  14'h024a;
         mem[2255] = -14'h0099;
         mem[2256] =  14'h005f;
         mem[2257] =  14'h000c;
         mem[2258] = -14'h0012;
         mem[2259] = -14'h000b;
         mem[2260] = -14'h00cc;
         mem[2261] = -14'h00a1;
         mem[2262] = -14'h000a;
         mem[2263] = -14'h0194;
         mem[2264] = -14'h000c;
         mem[2265] = -14'h0008;
         mem[2266] =  14'h002b;
         mem[2267] =  14'h0029;
         mem[2268] =  14'h0090;
         mem[2269] =  14'h001e;
         mem[2270] =  14'h00ed;
         mem[2271] = -14'h0029;
         mem[2272] =  14'h0104;
         mem[2273] =  14'h0008;
         mem[2274] = -14'h0002;
         mem[2275] = -14'h001d;
         mem[2276] = -14'h0011;
         mem[2277] = -14'h00ac;
         mem[2278] = -14'h00be;
         mem[2279] = -14'h0006;
         mem[2280] = -14'h0036;
         mem[2281] =  14'h0024;
         mem[2282] = -14'h0011;
         mem[2283] = -14'h0243;
         mem[2284] = -14'h0026;
         mem[2285] =  14'h006a;
         mem[2286] = -14'h006a;
         mem[2287] =  14'h000f;
         mem[2288] =  14'h0076;
         mem[2289] = -14'h0152;
         mem[2290] =  14'h0031;
         mem[2291] =  14'h0013;
         mem[2292] =  14'h0075;
         mem[2293] = -14'h007f;
         mem[2294] = -14'h018a;
         mem[2295] =  14'h001d;
         mem[2296] = -14'h0177;
         mem[2297] = -14'h001c;
         mem[2298] =  14'h0092;
         mem[2299] =  14'h0018;
         mem[2300] =  14'h00de;
         mem[2301] =  14'h000e;
         mem[2302] = -14'h0047;
         mem[2303] =  14'h004b;
         mem[2304] =  14'h009b;
         mem[2305] =  14'h0064;
         mem[2306] =  14'h0096;
         mem[2307] =  14'h00a3;
         mem[2308] = -14'h0025;
         mem[2309] = -14'h004a;
         mem[2310] =  14'h0086;
         mem[2311] = -14'h00e4;
         mem[2312] =  14'h0071;
         mem[2313] =  14'h002d;
         mem[2314] = -14'h004c;
         mem[2315] =  14'h0199;
         mem[2316] = -14'h0088;
         mem[2317] = -14'h006b;
         mem[2318] =  14'h0021;
         mem[2319] =  14'h00fb;
         mem[2320] = -14'h0090;
         mem[2321] = -14'h0002;
         mem[2322] =  14'h0022;
         mem[2323] =  14'h0018;
         mem[2324] = -14'h000a;
         mem[2325] = -14'h0007;
         mem[2326] =  14'h0039;
         mem[2327] = -14'h0007;
         mem[2328] =  14'h0020;
         mem[2329] =  14'h0041;
         mem[2330] =  14'h0027;
         mem[2331] =  14'h0000;
         mem[2332] = -14'h008d;
         mem[2333] = -14'h002c;
         mem[2334] =  14'h000a;
         mem[2335] = -14'h0003;
         mem[2336] = -14'h0004;
         mem[2337] =  14'h0023;
         mem[2338] =  14'h003c;
         mem[2339] = -14'h014b;
         mem[2340] = -14'h002f;
         mem[2341] = -14'h0032;
         mem[2342] = -14'h0053;
         mem[2343] = -14'h0001;
         mem[2344] =  14'h0097;
         mem[2345] = -14'h003c;
         mem[2346] =  14'h00bb;
         mem[2347] =  14'h0117;
         mem[2348] =  14'h002b;
         mem[2349] =  14'h0101;
         mem[2350] = -14'h000d;
         mem[2351] = -14'h00f0;
         mem[2352] =  14'h008b;
         mem[2353] =  14'h0067;
         mem[2354] =  14'h0008;
         mem[2355] = -14'h0059;
         mem[2356] =  14'h002b;
         mem[2357] = -14'h0033;
         mem[2358] = -14'h007e;
         mem[2359] = -14'h0004;
         mem[2360] = -14'h002a;
         mem[2361] = -14'h006a;
         mem[2362] =  14'h00b5;
         mem[2363] = -14'h004e;
         mem[2364] =  14'h0006;
         mem[2365] = -14'h002a;
         mem[2366] =  14'h0033;
         mem[2367] =  14'h0001;
         mem[2368] =  14'h00e0;
         mem[2369] = -14'h002c;
         mem[2370] = -14'h009b;
         mem[2371] = -14'h0031;
         mem[2372] =  14'h0029;
         mem[2373] = -14'h00c4;
         mem[2374] = -14'h001d;
         mem[2375] = -14'h0009;
         mem[2376] =  14'h002f;
         mem[2377] =  14'h0001;
         mem[2378] =  14'h001f;
         mem[2379] = -14'h0031;
         mem[2380] =  14'h003e;
         mem[2381] = -14'h0063;
         mem[2382] = -14'h1e00;
         mem[2383] = -14'h0010;
         mem[2384] = -14'h00b3;
         mem[2385] =  14'h000f;
         mem[2386] =  14'h0000;
         mem[2387] = -14'h0024;
         mem[2388] =  14'h0000;
         mem[2389] = -14'h0004;
         mem[2390] = -14'h006b;
         mem[2391] = -14'h0034;
         mem[2392] =  14'h002d;
         mem[2393] =  14'h0007;
         mem[2394] =  14'h004d;
         mem[2395] = -14'h0043;
         mem[2396] =  14'h0012;
         mem[2397] = -14'h00db;
         mem[2398] = -14'h000c;
         mem[2399] = -14'h0073;
         mem[2400] = -14'h0077;
         mem[2401] = -14'h000b;
         mem[2402] =  14'h0049;
         mem[2403] = -14'h0002;
         mem[2404] = -14'h0386;
         mem[2405] =  14'h0177;
         mem[2406] = -14'h014d;
         mem[2407] = -14'h0002;
         mem[2408] =  14'h0015;
         mem[2409] = -14'h002b;
         mem[2410] =  14'h0040;
         mem[2411] = -14'h003e;
         mem[2412] =  14'h0033;
         mem[2413] = -14'h0110;
         mem[2414] =  14'h007f;
         mem[2415] =  14'h006a;
         mem[2416] =  14'h0022;
         mem[2417] =  14'h0095;
         mem[2418] = -14'h0325;
         mem[2419] =  14'h00b1;
         mem[2420] =  14'h004d;
         mem[2421] = -14'h0051;
         mem[2422] =  14'h000e;
         mem[2423] =  14'h00eb;
         mem[2424] =  14'h0033;
         mem[2425] =  14'h0005;
         mem[2426] =  14'h0021;
         mem[2427] = -14'h0031;
         mem[2428] =  14'h0028;
         mem[2429] = -14'h008d;
         mem[2430] = -14'h000b;
         mem[2431] = -14'h00f1;
         mem[2432] = -14'h0001;
         mem[2433] = -14'h0005;
         mem[2434] =  14'h001c;
         mem[2435] =  14'h0002;
         mem[2436] = -14'h0015;
         mem[2437] =  14'h0122;
         mem[2438] =  14'h00c3;
         mem[2439] = -14'h000f;
         mem[2440] =  14'h0017;
         mem[2441] =  14'h0015;
         mem[2442] = -14'h0119;
         mem[2443] = -14'h0033;
         mem[2444] =  14'h0024;
         mem[2445] = -14'h013b;
         mem[2446] =  14'h0003;
         mem[2447] = -14'h0052;
         mem[2448] =  14'h003a;
         mem[2449] =  14'h0082;
         mem[2450] =  14'h0012;
         mem[2451] =  14'h0028;
         mem[2452] = -14'h002d;
         mem[2453] =  14'h000e;
         mem[2454] = -14'h0012;
         mem[2455] = -14'h0032;
         mem[2456] = -14'h00dc;
         mem[2457] = -14'h0122;
         mem[2458] =  14'h0028;
         mem[2459] = -14'h009d;
         mem[2460] =  14'h00b2;
         mem[2461] = -14'h0026;
         mem[2462] =  14'h002c;
         mem[2463] =  14'h009e;
         mem[2464] =  14'h006c;
         mem[2465] =  14'h0140;
         mem[2466] =  14'h0024;
         mem[2467] =  14'h0098;
         mem[2468] = -14'h00c9;
         mem[2469] = -14'h016c;
         mem[2470] =  14'h0007;
         mem[2471] = -14'h0039;
         mem[2472] =  14'h0051;
         mem[2473] =  14'h00a6;
         mem[2474] =  14'h001c;
         mem[2475] =  14'h0005;
         mem[2476] =  14'h0008;
         mem[2477] = -14'h0041;
         mem[2478] =  14'h00e8;
         mem[2479] =  14'h0002;
         mem[2480] = -14'h00f5;
         mem[2481] =  14'h015e;
         mem[2482] =  14'h0037;
         mem[2483] = -14'h00e2;
         mem[2484] =  14'h0010;
         mem[2485] = -14'h0026;
         mem[2486] =  14'h0020;
         mem[2487] = -14'h0010;
         mem[2488] =  14'h001c;
         mem[2489] =  14'h005d;
         mem[2490] =  14'h0046;
         mem[2491] =  14'h0114;
         mem[2492] =  14'h0034;
         mem[2493] =  14'h0006;
         mem[2494] =  14'h000e;
         mem[2495] =  14'h0035;
         mem[2496] = -14'h0190;
         mem[2497] =  14'h0086;
         mem[2498] = -14'h014f;
         mem[2499] = -14'h0082;
         mem[2500] =  14'h0010;
         mem[2501] =  14'h0313;
         mem[2502] =  14'h0063;
         mem[2503] =  14'h0073;
         mem[2504] =  14'h006d;
         mem[2505] = -14'h00aa;
         mem[2506] =  14'h0047;
         mem[2507] =  14'h0071;
         mem[2508] = -14'h0040;
         mem[2509] =  14'h0058;
         mem[2510] =  14'h0008;
         mem[2511] = -14'h000f;
         mem[2512] = -14'h003e;
         mem[2513] = -14'h007b;
         mem[2514] =  14'h00b8;
         mem[2515] = -14'h0057;
         mem[2516] = -14'h00d2;
         mem[2517] =  14'h0030;
         mem[2518] = -14'h0007;
         mem[2519] = -14'h008a;
         mem[2520] = -14'h000a;
         mem[2521] =  14'h0027;
         mem[2522] = -14'h0038;
         mem[2523] =  14'h009b;
         mem[2524] = -14'h0003;
         mem[2525] = -14'h0046;
         mem[2526] = -14'h000a;
         mem[2527] = -14'h000e;
         mem[2528] = -14'h008c;
         mem[2529] =  14'h007b;
         mem[2530] = -14'h0054;
         mem[2531] =  14'h0020;
         mem[2532] =  14'h008a;
         mem[2533] =  14'h000b;
         mem[2534] =  14'h006a;
         mem[2535] =  14'h00b0;
         mem[2536] = -14'h003a;
         mem[2537] = -14'h0037;
         mem[2538] = -14'h00b9;
         mem[2539] =  14'h002f;
         mem[2540] = -14'h0076;
         mem[2541] =  14'h003d;
         mem[2542] =  14'h0008;
         mem[2543] =  14'h0013;
         mem[2544] = -14'h002f;
         mem[2545] = -14'h1e00;
         mem[2546] = -14'h000c;
         mem[2547] =  14'h0028;
         mem[2548] = -14'h0040;
         mem[2549] =  14'h002f;
         mem[2550] = -14'h0031;
         mem[2551] =  14'h003a;
         mem[2552] = -14'h00aa;
         mem[2553] =  14'h00a5;
         mem[2554] =  14'h0059;
         mem[2555] =  14'h0035;
         mem[2556] = -14'h002d;
         mem[2557] =  14'h004e;
         mem[2558] =  14'h0100;
         mem[2559] = -14'h0010;
         mem[2560] = -14'h004e;
         mem[2561] = -14'h00f0;
         mem[2562] = -14'h0006;
         mem[2563] =  14'h0015;
         mem[2564] = -14'h004f;
         mem[2565] = -14'h00d8;
         mem[2566] = -14'h0156;
         mem[2567] = -14'h009b;
         mem[2568] = -14'h0009;
         mem[2569] =  14'h0053;
         mem[2570] =  14'h004b;
         mem[2571] = -14'h0180;
         mem[2572] = -14'h000b;
         mem[2573] = -14'h0025;
         mem[2574] = -14'h0009;
         mem[2575] =  14'h0099;
         mem[2576] = -14'h0009;
         mem[2577] =  14'h000e;
         mem[2578] = -14'h0043;
         mem[2579] =  14'h005b;
         mem[2580] =  14'h0083;
         mem[2581] =  14'h0000;
         mem[2582] =  14'h009d;
         mem[2583] =  14'h002e;
         mem[2584] = -14'h01ed;
         mem[2585] =  14'h009d;
         mem[2586] =  14'h0071;
         mem[2587] =  14'h003e;
         mem[2588] = -14'h0026;
         mem[2589] = -14'h002e;
         mem[2590] = -14'h0030;
         mem[2591] =  14'h003a;
         mem[2592] = -14'h0084;
         mem[2593] =  14'h0059;
         mem[2594] = -14'h0037;
         mem[2595] = -14'h0049;
         mem[2596] =  14'h0043;
         mem[2597] = -14'h007f;
         mem[2598] = -14'h00c5;
         mem[2599] = -14'h0052;
         mem[2600] = -14'h0039;
         mem[2601] =  14'h0083;
         mem[2602] =  14'h000c;
         mem[2603] =  14'h0001;
         mem[2604] =  14'h0011;
         mem[2605] = -14'h01e5;
         mem[2606] = -14'h016d;
         mem[2607] =  14'h002e;
         mem[2608] = -14'h002a;
         mem[2609] = -14'h0047;
         mem[2610] = -14'h0004;
         mem[2611] = -14'h0001;
         mem[2612] =  14'h028a;
         mem[2613] =  14'h0049;
         mem[2614] =  14'h00a7;
         mem[2615] =  14'h0045;
         mem[2616] = -14'h0040;
         mem[2617] =  14'h000e;
         mem[2618] =  14'h0077;
         mem[2619] =  14'h0041;
         mem[2620] =  14'h0012;
         mem[2621] =  14'h002b;
         mem[2622] = -14'h002d;
         mem[2623] =  14'h0263;
         mem[2624] =  14'h009f;
         mem[2625] = -14'h0010;
         mem[2626] =  14'h001b;
         mem[2627] = -14'h00ea;
         mem[2628] =  14'h017d;
         mem[2629] =  14'h0032;
         mem[2630] =  14'h0000;
         mem[2631] =  14'h010b;
         mem[2632] =  14'h0045;
         mem[2633] =  14'h000e;
         mem[2634] = -14'h00f7;
         mem[2635] = -14'h0059;
         mem[2636] = -14'h000d;
         mem[2637] =  14'h0047;
         mem[2638] =  14'h0035;
         mem[2639] =  14'h001d;
         mem[2640] = -14'h0039;
         mem[2641] = -14'h0019;
         mem[2642] =  14'h0014;
         mem[2643] =  14'h0029;
         mem[2644] = -14'h002c;
         mem[2645] =  14'h0020;
         mem[2646] = -14'h011c;
         mem[2647] = -14'h04d2;
         mem[2648] = -14'h00a3;
         mem[2649] =  14'h0274;
         mem[2650] = -14'h0082;
         mem[2651] =  14'h001c;
         mem[2652] = -14'h016a;
         mem[2653] =  14'h000a;
         mem[2654] =  14'h0055;
         mem[2655] =  14'h000b;
         mem[2656] =  14'h0000;
         mem[2657] =  14'h005b;
         mem[2658] =  14'h0070;
         mem[2659] = -14'h000b;
         mem[2660] = -14'h00eb;
         mem[2661] =  14'h0033;
         mem[2662] = -14'h003b;
         mem[2663] =  14'h0044;
         mem[2664] =  14'h000c;
         mem[2665] = -14'h02d4;
         mem[2666] = -14'h0028;
         mem[2667] = -14'h01fe;
         mem[2668] =  14'h014e;
         mem[2669] = -14'h000b;
         mem[2670] = -14'h0034;
         mem[2671] = -14'h00f4;
         mem[2672] = -14'h021d;
         mem[2673] = -14'h019c;
         mem[2674] =  14'h00b3;
         mem[2675] = -14'h0066;
         mem[2676] =  14'h0071;
         mem[2677] = -14'h0193;
         mem[2678] = -14'h000a;
         mem[2679] = -14'h0003;
         mem[2680] =  14'h0006;
         mem[2681] = -14'h0010;
         mem[2682] = -14'h00d7;
         mem[2683] =  14'h0029;
         mem[2684] =  14'h0001;
         mem[2685] =  14'h0022;
         mem[2686] = -14'h0029;
         mem[2687] =  14'h008d;
         mem[2688] = -14'h0113;
         mem[2689] =  14'h012b;
         mem[2690] =  14'h0061;
         mem[2691] =  14'h001c;
         mem[2692] = -14'h002f;
         mem[2693] =  14'h002f;
         mem[2694] =  14'h00f3;
         mem[2695] =  14'h0009;
         mem[2696] = -14'h0010;
         mem[2697] =  14'h006b;
         mem[2698] = -14'h0036;
         mem[2699] = -14'h0220;
         mem[2700] = -14'h017c;
         mem[2701] =  14'h0052;
         mem[2702] =  14'h0030;
         mem[2703] =  14'h0047;
         mem[2704] =  14'h0044;
         mem[2705] = -14'h009b;
         mem[2706] =  14'h0005;
         mem[2707] =  14'h007c;
         mem[2708] = -14'h00ee;
         mem[2709] =  14'h0057;
         mem[2710] = -14'h000f;
         mem[2711] =  14'h00a4;
         mem[2712] = -14'h0065;
         mem[2713] = -14'h0075;
         mem[2714] =  14'h0037;
         mem[2715] =  14'h006c;
         mem[2716] = -14'h00a2;
         mem[2717] = -14'h004d;
         mem[2718] =  14'h0067;
         mem[2719] = -14'h00c7;
         mem[2720] =  14'h0029;
         mem[2721] = -14'h00cc;
         mem[2722] =  14'h0041;
         mem[2723] = -14'h00b5;
         mem[2724] =  14'h00bd;
         mem[2725] = -14'h003e;
         mem[2726] = -14'h0021;
         mem[2727] =  14'h0023;
         mem[2728] =  14'h00e5;
         mem[2729] = -14'h00dc;
         mem[2730] =  14'h00da;
         mem[2731] = -14'h004b;
         mem[2732] =  14'h0031;
         mem[2733] = -14'h0041;
         mem[2734] =  14'h0037;
         mem[2735] = -14'h000b;
         mem[2736] =  14'h0030;
         mem[2737] =  14'h0050;
         mem[2738] =  14'h002a;
         mem[2739] = -14'h009f;
         mem[2740] =  14'h0031;
         mem[2741] = -14'h0003;
         mem[2742] = -14'h0008;
         mem[2743] =  14'h0035;
         mem[2744] =  14'h002f;
         mem[2745] =  14'h000d;
         mem[2746] =  14'h0031;
         mem[2747] =  14'h00f4;
         mem[2748] =  14'h003f;
         mem[2749] = -14'h01a3;
         mem[2750] = -14'h0017;
         mem[2751] = -14'h005b;
         mem[2752] =  14'h0033;
         mem[2753] = -14'h0030;
         mem[2754] =  14'h00d1;
         mem[2755] = -14'h0075;
         mem[2756] =  14'h0024;
         mem[2757] = -14'h0034;
         mem[2758] =  14'h000d;
         mem[2759] = -14'h0038;
         mem[2760] =  14'h0024;
         mem[2761] =  14'h01ca;
         mem[2762] = -14'h01e3;
         mem[2763] = -14'h000e;
         mem[2764] = -14'h001a;
         mem[2765] = -14'h000c;
         mem[2766] = -14'h0017;
         mem[2767] = -14'h016d;
         mem[2768] =  14'h0052;
         mem[2769] = -14'h0008;
         mem[2770] = -14'h0004;
         mem[2771] =  14'h0117;
         mem[2772] =  14'h004f;
         mem[2773] = -14'h00b0;
         mem[2774] = -14'h0001;
         mem[2775] =  14'h0020;
         mem[2776] =  14'h0064;
         mem[2777] = -14'h0033;
         mem[2778] =  14'h00e8;
         mem[2779] = -14'h0032;
         mem[2780] = -14'h0084;
         mem[2781] = -14'h0008;
         mem[2782] =  14'h0020;
         mem[2783] = -14'h00a2;
         mem[2784] =  14'h0010;
         mem[2785] =  14'h004f;
         mem[2786] =  14'h002b;
         mem[2787] =  14'h005a;
         mem[2788] = -14'h00be;
         mem[2789] =  14'h006a;
         mem[2790] =  14'h0000;
         mem[2791] = -14'h002a;
         mem[2792] = -14'h0085;
         mem[2793] =  14'h0000;
         mem[2794] =  14'h000f;
         mem[2795] =  14'h0025;
         mem[2796] =  14'h0021;
         mem[2797] = -14'h015e;
         mem[2798] = -14'h0001;
         mem[2799] = -14'h004f;
         mem[2800] =  14'h0015;
         mem[2801] = -14'h002d;
         mem[2802] =  14'h0024;
         mem[2803] = -14'h003c;
         mem[2804] = -14'h0005;
         mem[2805] = -14'h0005;
         mem[2806] =  14'h0076;
         mem[2807] =  14'h0066;
         mem[2808] =  14'h0007;
         mem[2809] =  14'h006f;
         mem[2810] =  14'h0011;
         mem[2811] = -14'h0035;
         mem[2812] =  14'h005c;
         mem[2813] = -14'h0027;
         mem[2814] =  14'h0047;
         mem[2815] = -14'h005d;
         mem[2816] =  14'h006a;
         mem[2817] = -14'h002b;
         mem[2818] = -14'h00a7;
         mem[2819] = -14'h0075;
         mem[2820] =  14'h0012;
         mem[2821] = -14'h0101;
         mem[2822] =  14'h006c;
         mem[2823] =  14'h0043;
         mem[2824] = -14'h010a;
         mem[2825] = -14'h0005;
         mem[2826] =  14'h0190;
         mem[2827] =  14'h0025;
         mem[2828] =  14'h0000;
         mem[2829] = -14'h0009;
         mem[2830] = -14'h00df;
         mem[2831] =  14'h0098;
         mem[2832] = -14'h000e;
         mem[2833] = -14'h015c;
         mem[2834] =  14'h0041;
         mem[2835] = -14'h0024;
         mem[2836] =  14'h002b;
         mem[2837] =  14'h0049;
         mem[2838] =  14'h0034;
         mem[2839] = -14'h0027;
         mem[2840] =  14'h0013;
         mem[2841] =  14'h0014;
         mem[2842] = -14'h005e;
         mem[2843] = -14'h00ec;
         mem[2844] =  14'h0014;
         mem[2845] =  14'h00b7;
         mem[2846] = -14'h00e0;
         mem[2847] = -14'h0097;
         mem[2848] =  14'h007b;
         mem[2849] =  14'h0056;
         mem[2850] =  14'h0050;
         mem[2851] =  14'h002d;
         mem[2852] = -14'h004b;
         mem[2853] = -14'h0024;
         mem[2854] =  14'h008e;
         mem[2855] = -14'h0010;
         mem[2856] =  14'h0032;
         mem[2857] =  14'h004b;
         mem[2858] =  14'h00ab;
         mem[2859] =  14'h0000;
         mem[2860] =  14'h001e;
         mem[2861] = -14'h0081;
         mem[2862] = -14'h0037;
         mem[2863] = -14'h0026;
         mem[2864] =  14'h0066;
         mem[2865] =  14'h001d;
         mem[2866] =  14'h0015;
         mem[2867] = -14'h0030;
         mem[2868] =  14'h0028;
         mem[2869] = -14'h0111;
         mem[2870] =  14'h000d;
         mem[2871] = -14'h000f;
         mem[2872] =  14'h00a9;
         mem[2873] =  14'h000f;
         mem[2874] = -14'h003f;
         mem[2875] =  14'h0065;
         mem[2876] = -14'h0018;
         mem[2877] = -14'h0075;
         mem[2878] =  14'h0025;
         mem[2879] =  14'h0194;
         mem[2880] =  14'h0013;
         mem[2881] =  14'h0078;
         mem[2882] =  14'h001e;
         mem[2883] = -14'h00d6;
         mem[2884] =  14'h0014;
         mem[2885] = -14'h002d;
         mem[2886] =  14'h0020;
         mem[2887] =  14'h0045;
         mem[2888] = -14'h006e;
         mem[2889] =  14'h0096;
         mem[2890] = -14'h0009;
         mem[2891] = -14'h0005;
         mem[2892] =  14'h0024;
         mem[2893] = -14'h006a;
         mem[2894] =  14'h0035;
         mem[2895] =  14'h00a2;
         mem[2896] = -14'h0083;
         mem[2897] = -14'h002d;
         mem[2898] =  14'h00af;
         mem[2899] = -14'h0028;
         mem[2900] = -14'h003e;
         mem[2901] = -14'h00e1;
         mem[2902] =  14'h002d;
         mem[2903] = -14'h002a;
         mem[2904] =  14'h0058;
         mem[2905] =  14'h00dd;
         mem[2906] =  14'h001e;
         mem[2907] = -14'h00e6;
         mem[2908] = -14'h0115;
         mem[2909] = -14'h0008;
         mem[2910] =  14'h0037;
         mem[2911] =  14'h01ae;
         mem[2912] =  14'h0000;
     end

endmodule: leafVal0_rom
