module rect0_rom
  #(
     parameter W_DATA = 5,
     parameter W_ADDR = 14
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1

     );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               14'b00000000000000: data1 <= 5'h06;
               14'b00000000000001: data1 <= 5'h04;
               14'b00000000000010: data1 <= 5'h0c;
               14'b00000000000011: data1 <= 5'h09;
               14'b00000000000100: data1 <= 5'h06;
               14'b00000000000101: data1 <= 5'h04;
               14'b00000000000110: data1 <= 5'h0c;
               14'b00000000000111: data1 <= 5'h07;
               14'b00000000001000: data1 <= 5'h03;
               14'b00000000001001: data1 <= 5'h09;
               14'b00000000001010: data1 <= 5'h12;
               14'b00000000001011: data1 <= 5'h09;
               14'b00000000001100: data1 <= 5'h08;
               14'b00000000001101: data1 <= 5'h12;
               14'b00000000001110: data1 <= 5'h09;
               14'b00000000001111: data1 <= 5'h06;
               14'b00000000010000: data1 <= 5'h03;
               14'b00000000010001: data1 <= 5'h05;
               14'b00000000010010: data1 <= 5'h04;
               14'b00000000010011: data1 <= 5'h13;
               14'b00000000010100: data1 <= 5'h06;
               14'b00000000010101: data1 <= 5'h05;
               14'b00000000010110: data1 <= 5'h0c;
               14'b00000000010111: data1 <= 5'h10;
               14'b00000000011000: data1 <= 5'h05;
               14'b00000000011001: data1 <= 5'h08;
               14'b00000000011010: data1 <= 5'h0c;
               14'b00000000011011: data1 <= 5'h06;
               14'b00000000011100: data1 <= 5'h0b;
               14'b00000000011101: data1 <= 5'h0e;
               14'b00000000011110: data1 <= 5'h04;
               14'b00000000011111: data1 <= 5'h0a;
               14'b00000000100000: data1 <= 5'h04;
               14'b00000000100001: data1 <= 5'h00;
               14'b00000000100010: data1 <= 5'h07;
               14'b00000000100011: data1 <= 5'h06;
               14'b00000000100100: data1 <= 5'h06;
               14'b00000000100101: data1 <= 5'h06;
               14'b00000000100110: data1 <= 5'h0c;
               14'b00000000100111: data1 <= 5'h06;
               14'b00000000101000: data1 <= 5'h06;
               14'b00000000101001: data1 <= 5'h04;
               14'b00000000101010: data1 <= 5'h0c;
               14'b00000000101011: data1 <= 5'h07;
               14'b00000000101100: data1 <= 5'h01;
               14'b00000000101101: data1 <= 5'h08;
               14'b00000000101110: data1 <= 5'h13;
               14'b00000000101111: data1 <= 5'h0c;
               14'b00000000110000: data1 <= 5'h00;
               14'b00000000110001: data1 <= 5'h02;
               14'b00000000110010: data1 <= 5'h18;
               14'b00000000110011: data1 <= 5'h03;
               14'b00000000110100: data1 <= 5'h09;
               14'b00000000110101: data1 <= 5'h09;
               14'b00000000110110: data1 <= 5'h06;
               14'b00000000110111: data1 <= 5'h0f;
               14'b00000000111000: data1 <= 5'h05;
               14'b00000000111001: data1 <= 5'h06;
               14'b00000000111010: data1 <= 5'h0e;
               14'b00000000111011: data1 <= 5'h0a;
               14'b00000000111100: data1 <= 5'h05;
               14'b00000000111101: data1 <= 5'h00;
               14'b00000000111110: data1 <= 5'h0e;
               14'b00000000111111: data1 <= 5'h09;
               14'b00000001000000: data1 <= 5'h0d;
               14'b00000001000001: data1 <= 5'h0b;
               14'b00000001000010: data1 <= 5'h09;
               14'b00000001000011: data1 <= 5'h06;
               14'b00000001000100: data1 <= 5'h07;
               14'b00000001000101: data1 <= 5'h05;
               14'b00000001000110: data1 <= 5'h06;
               14'b00000001000111: data1 <= 5'h0a;
               14'b00000001001000: data1 <= 5'h0a;
               14'b00000001001001: data1 <= 5'h08;
               14'b00000001001010: data1 <= 5'h06;
               14'b00000001001011: data1 <= 5'h0a;
               14'b00000001001100: data1 <= 5'h02;
               14'b00000001001101: data1 <= 5'h05;
               14'b00000001001110: data1 <= 5'h04;
               14'b00000001001111: data1 <= 5'h09;
               14'b00000001010000: data1 <= 5'h12;
               14'b00000001010001: data1 <= 5'h00;
               14'b00000001010010: data1 <= 5'h06;
               14'b00000001010011: data1 <= 5'h0b;
               14'b00000001010100: data1 <= 5'h00;
               14'b00000001010101: data1 <= 5'h06;
               14'b00000001010110: data1 <= 5'h18;
               14'b00000001010111: data1 <= 5'h0d;
               14'b00000001011000: data1 <= 5'h09;
               14'b00000001011001: data1 <= 5'h06;
               14'b00000001011010: data1 <= 5'h06;
               14'b00000001011011: data1 <= 5'h09;
               14'b00000001011100: data1 <= 5'h07;
               14'b00000001011101: data1 <= 5'h12;
               14'b00000001011110: data1 <= 5'h0a;
               14'b00000001011111: data1 <= 5'h06;
               14'b00000001100000: data1 <= 5'h05;
               14'b00000001100001: data1 <= 5'h07;
               14'b00000001100010: data1 <= 5'h0e;
               14'b00000001100011: data1 <= 5'h0c;
               14'b00000001100100: data1 <= 5'h00;
               14'b00000001100101: data1 <= 5'h03;
               14'b00000001100110: data1 <= 5'h18;
               14'b00000001100111: data1 <= 5'h03;
               14'b00000001101000: data1 <= 5'h05;
               14'b00000001101001: data1 <= 5'h08;
               14'b00000001101010: data1 <= 5'h0f;
               14'b00000001101011: data1 <= 5'h06;
               14'b00000001101100: data1 <= 5'h09;
               14'b00000001101101: data1 <= 5'h06;
               14'b00000001101110: data1 <= 5'h05;
               14'b00000001101111: data1 <= 5'h0e;
               14'b00000001110000: data1 <= 5'h09;
               14'b00000001110001: data1 <= 5'h05;
               14'b00000001110010: data1 <= 5'h06;
               14'b00000001110011: data1 <= 5'h0a;
               14'b00000001110100: data1 <= 5'h06;
               14'b00000001110101: data1 <= 5'h06;
               14'b00000001110110: data1 <= 5'h03;
               14'b00000001110111: data1 <= 5'h0c;
               14'b00000001111000: data1 <= 5'h03;
               14'b00000001111001: data1 <= 5'h15;
               14'b00000001111010: data1 <= 5'h12;
               14'b00000001111011: data1 <= 5'h03;
               14'b00000001111100: data1 <= 5'h05;
               14'b00000001111101: data1 <= 5'h06;
               14'b00000001111110: data1 <= 5'h0d;
               14'b00000001111111: data1 <= 5'h06;
               14'b00000010000000: data1 <= 5'h12;
               14'b00000010000001: data1 <= 5'h01;
               14'b00000010000010: data1 <= 5'h06;
               14'b00000010000011: data1 <= 5'h0f;
               14'b00000010000100: data1 <= 5'h01;
               14'b00000010000101: data1 <= 5'h01;
               14'b00000010000110: data1 <= 5'h06;
               14'b00000010000111: data1 <= 5'h0f;
               14'b00000010001000: data1 <= 5'h00;
               14'b00000010001001: data1 <= 5'h08;
               14'b00000010001010: data1 <= 5'h18;
               14'b00000010001011: data1 <= 5'h0f;
               14'b00000010001100: data1 <= 5'h05;
               14'b00000010001101: data1 <= 5'h06;
               14'b00000010001110: data1 <= 5'h0e;
               14'b00000010001111: data1 <= 5'h0c;
               14'b00000010010000: data1 <= 5'h02;
               14'b00000010010001: data1 <= 5'h0c;
               14'b00000010010010: data1 <= 5'h15;
               14'b00000010010011: data1 <= 5'h0c;
               14'b00000010010100: data1 <= 5'h08;
               14'b00000010010101: data1 <= 5'h01;
               14'b00000010010110: data1 <= 5'h04;
               14'b00000010010111: data1 <= 5'h0a;
               14'b00000010011000: data1 <= 5'h02;
               14'b00000010011001: data1 <= 5'h0d;
               14'b00000010011010: data1 <= 5'h14;
               14'b00000010011011: data1 <= 5'h0a;
               14'b00000010011100: data1 <= 5'h00;
               14'b00000010011101: data1 <= 5'h01;
               14'b00000010011110: data1 <= 5'h06;
               14'b00000010011111: data1 <= 5'h0d;
               14'b00000010100000: data1 <= 5'h14;
               14'b00000010100001: data1 <= 5'h02;
               14'b00000010100010: data1 <= 5'h04;
               14'b00000010100011: data1 <= 5'h0d;
               14'b00000010100100: data1 <= 5'h00;
               14'b00000010100101: data1 <= 5'h05;
               14'b00000010100110: data1 <= 5'h16;
               14'b00000010100111: data1 <= 5'h13;
               14'b00000010101000: data1 <= 5'h12;
               14'b00000010101001: data1 <= 5'h04;
               14'b00000010101010: data1 <= 5'h06;
               14'b00000010101011: data1 <= 5'h09;
               14'b00000010101100: data1 <= 5'h00;
               14'b00000010101101: data1 <= 5'h03;
               14'b00000010101110: data1 <= 5'h06;
               14'b00000010101111: data1 <= 5'h0b;
               14'b00000010110000: data1 <= 5'h0c;
               14'b00000010110001: data1 <= 5'h01;
               14'b00000010110010: data1 <= 5'h04;
               14'b00000010110011: data1 <= 5'h09;
               14'b00000010110100: data1 <= 5'h00;
               14'b00000010110101: data1 <= 5'h06;
               14'b00000010110110: data1 <= 5'h13;
               14'b00000010110111: data1 <= 5'h03;
               14'b00000010111000: data1 <= 5'h0c;
               14'b00000010111001: data1 <= 5'h01;
               14'b00000010111010: data1 <= 5'h04;
               14'b00000010111011: data1 <= 5'h09;
               14'b00000010111100: data1 <= 5'h08;
               14'b00000010111101: data1 <= 5'h01;
               14'b00000010111110: data1 <= 5'h04;
               14'b00000010111111: data1 <= 5'h09;
               14'b00000011000000: data1 <= 5'h05;
               14'b00000011000001: data1 <= 5'h05;
               14'b00000011000010: data1 <= 5'h0e;
               14'b00000011000011: data1 <= 5'h0e;
               14'b00000011000100: data1 <= 5'h01;
               14'b00000011000101: data1 <= 5'h0a;
               14'b00000011000110: data1 <= 5'h12;
               14'b00000011000111: data1 <= 5'h02;
               14'b00000011001000: data1 <= 5'h11;
               14'b00000011001001: data1 <= 5'h0d;
               14'b00000011001010: data1 <= 5'h04;
               14'b00000011001011: data1 <= 5'h0b;
               14'b00000011001100: data1 <= 5'h00;
               14'b00000011001101: data1 <= 5'h04;
               14'b00000011001110: data1 <= 5'h06;
               14'b00000011001111: data1 <= 5'h09;
               default: data1 <= 0;
           endcase
        end

endmodule: rect0_rom
