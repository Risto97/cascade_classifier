module leafVal0_rom
  #(
     parameter W_DATA = 11,
     parameter W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               8'b00000000: data1 <= -11'h237;
               8'b00000001: data1 <=  11'h153;
               8'b00000010: data1 <=  11'h110;
               8'b00000011: data1 <=  11'h12d;
               8'b00000100: data1 <=  11'h142;
               8'b00000101: data1 <= -11'h1df;
               8'b00000110: data1 <=  11'h070;
               8'b00000111: data1 <=  11'h071;
               8'b00001000: data1 <=  11'h0da;
               8'b00001001: data1 <= -11'h192;
               8'b00001010: data1 <=  11'h12e;
               8'b00001011: data1 <=  11'h0b3;
               8'b00001100: data1 <=  11'h1ba;
               8'b00001101: data1 <= -11'h22e;
               8'b00001110: data1 <=  11'h074;
               8'b00001111: data1 <=  11'h089;
               8'b00010000: data1 <=  11'h0ee;
               8'b00010001: data1 <= -11'h0a9;
               8'b00010010: data1 <= -11'h04c;
               8'b00010011: data1 <=  11'h15b;
               8'b00010100: data1 <= -11'h032;
               8'b00010101: data1 <= -11'h087;
               8'b00010110: data1 <=  11'h124;
               8'b00010111: data1 <=  11'h0c5;
               8'b00011000: data1 <= -11'h183;
               8'b00011001: data1 <=  11'h177;
               8'b00011010: data1 <=  11'h100;
               8'b00011011: data1 <= -11'h198;
               8'b00011100: data1 <=  11'h0d4;
               8'b00011101: data1 <=  11'h06c;
               8'b00011110: data1 <=  11'h10d;
               8'b00011111: data1 <= -11'h158;
               8'b00100000: data1 <=  11'h173;
               8'b00100001: data1 <=  11'h136;
               8'b00100010: data1 <= -11'h075;
               8'b00100011: data1 <=  11'h027;
               8'b00100100: data1 <= -11'h190;
               8'b00100101: data1 <=  11'h03b;
               8'b00100110: data1 <=  11'h147;
               8'b00100111: data1 <= -11'h04d;
               8'b00101000: data1 <= -11'h00d;
               8'b00101001: data1 <=  11'h189;
               8'b00101010: data1 <=  11'h0ef;
               8'b00101011: data1 <=  11'h0f6;
               8'b00101100: data1 <= -11'h2f5;
               8'b00101101: data1 <= -11'h070;
               8'b00101110: data1 <=  11'h066;
               8'b00101111: data1 <= -11'h2a5;
               8'b00110000: data1 <=  11'h048;
               8'b00110001: data1 <=  11'h03b;
               8'b00110010: data1 <=  11'h113;
               8'b00110011: data1 <=  11'h019;
               8'b00110100: data1 <= -11'h112;
               8'b00110101: data1 <=  11'h0c4;
               8'b00110110: data1 <=  11'h161;
               8'b00110111: data1 <=  11'h084;
               8'b00111000: data1 <=  11'h095;
               8'b00111001: data1 <=  11'h12b;
               8'b00111010: data1 <=  11'h0f4;
               8'b00111011: data1 <= -11'h023;
               8'b00111100: data1 <=  11'h046;
               8'b00111101: data1 <=  11'h03c;
               8'b00111110: data1 <= -11'h157;
               8'b00111111: data1 <= -11'h0e6;
               8'b01000000: data1 <= -11'h1a2;
               8'b01000001: data1 <=  11'h02e;
               8'b01000010: data1 <= -11'h061;
               8'b01000011: data1 <=  11'h03f;
               8'b01000100: data1 <= -11'h04b;
               8'b01000101: data1 <=  11'h0a1;
               8'b01000110: data1 <=  11'h00d;
               8'b01000111: data1 <=  11'h063;
               8'b01001000: data1 <=  11'h019;
               8'b01001001: data1 <= -11'h142;
               8'b01001010: data1 <= -11'h261;
               8'b01001011: data1 <= -11'h046;
               8'b01001100: data1 <= -11'h123;
               8'b01001101: data1 <= -11'h144;
               8'b01001110: data1 <=  11'h045;
               8'b01001111: data1 <=  11'h0b5;
               8'b01010000: data1 <=  11'h009;
               8'b01010001: data1 <= -11'h00c;
               8'b01010010: data1 <= -11'h059;
               8'b01010011: data1 <=  11'h036;
               8'b01010100: data1 <=  11'h115;
               8'b01010101: data1 <=  11'h167;
               8'b01010110: data1 <=  11'h0bd;
               8'b01010111: data1 <=  11'h060;
               8'b01011000: data1 <=  11'h143;
               8'b01011001: data1 <=  11'h075;
               8'b01011010: data1 <= -11'h0f5;
               8'b01011011: data1 <=  11'h00b;
               8'b01011100: data1 <=  11'h08a;
               8'b01011101: data1 <= -11'h17d;
               8'b01011110: data1 <= -11'h086;
               8'b01011111: data1 <= -11'h199;
               8'b01100000: data1 <=  11'h027;
               8'b01100001: data1 <= -11'h0b8;
               8'b01100010: data1 <=  11'h011;
               8'b01100011: data1 <=  11'h0ae;
               8'b01100100: data1 <=  11'h013;
               8'b01100101: data1 <= -11'h037;
               8'b01100110: data1 <=  11'h14f;
               8'b01100111: data1 <=  11'h138;
               8'b01101000: data1 <=  11'h0d9;
               8'b01101001: data1 <=  11'h04c;
               8'b01101010: data1 <= -11'h053;
               8'b01101011: data1 <= -11'h0d6;
               8'b01101100: data1 <= -11'h0ab;
               8'b01101101: data1 <=  11'h023;
               8'b01101110: data1 <=  11'h013;
               8'b01101111: data1 <=  11'h031;
               8'b01110000: data1 <=  11'h011;
               8'b01110001: data1 <=  11'h0c7;
               8'b01110010: data1 <=  11'h01f;
               8'b01110011: data1 <=  11'h003;
               8'b01110100: data1 <=  11'h087;
               8'b01110101: data1 <=  11'h064;
               8'b01110110: data1 <= -11'h21e;
               8'b01110111: data1 <=  11'h0fc;
               8'b01111000: data1 <=  11'h018;
               8'b01111001: data1 <= -11'h025;
               8'b01111010: data1 <= -11'h094;
               8'b01111011: data1 <= -11'h02b;
               8'b01111100: data1 <= -11'h0a3;
               8'b01111101: data1 <=  11'h040;
               8'b01111110: data1 <= -11'h045;
               8'b01111111: data1 <=  11'h03c;
               8'b10000000: data1 <= -11'h143;
               8'b10000001: data1 <=  11'h04d;
               8'b10000010: data1 <=  11'h087;
               8'b10000011: data1 <=  11'h03d;
               8'b10000100: data1 <=  11'h084;
               8'b10000101: data1 <= -11'h003;
               8'b10000110: data1 <= -11'h042;
               8'b10000111: data1 <= -11'h097;
               default: data1 <= 0;
           endcase
        end

endmodule: leafVal0_rom
