module featureThreshold_rom
  #(
     parameter W_DATA = 13,
     parameter W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1

     );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               12'b000000000000: data1 <= -13'h0081;
               12'b000000000001: data1 <= 13'h0032;
               12'b000000000010: data1 <= 13'h0059;
               12'b000000000011: data1 <= 13'h0017;
               12'b000000000100: data1 <= 13'h003d;
               12'b000000000101: data1 <= 13'h0197;
               12'b000000000110: data1 <= 13'h000b;
               12'b000000000111: data1 <= -13'h004d;
               12'b000000001000: data1 <= 13'h0018;
               12'b000000001001: data1 <= -13'h0056;
               12'b000000001010: data1 <= 13'h0053;
               12'b000000001011: data1 <= 13'h0057;
               12'b000000001100: data1 <= 13'h0177;
               12'b000000001101: data1 <= 13'h0094;
               12'b000000001110: data1 <= -13'h004e;
               12'b000000001111: data1 <= 13'h0021;
               12'b000000010000: data1 <= 13'h004b;
               12'b000000010001: data1 <= -13'h001c;
               12'b000000010010: data1 <= -13'h0028;
               12'b000000010011: data1 <= 13'h0040;
               12'b000000010100: data1 <= -13'h0054;
               12'b000000010101: data1 <= -13'h0233;
               12'b000000010110: data1 <= 13'h003a;
               12'b000000010111: data1 <= 13'h0029;
               12'b000000011000: data1 <= 13'h0176;
               12'b000000011001: data1 <= 13'h011d;
               12'b000000011010: data1 <= 13'h0081;
               12'b000000011011: data1 <= 13'h003a;
               12'b000000011100: data1 <= 13'h003b;
               12'b000000011101: data1 <= -13'h000c;
               12'b000000011110: data1 <= 13'h0086;
               12'b000000011111: data1 <= -13'h001d;
               12'b000000100000: data1 <= 13'h00ce;
               12'b000000100001: data1 <= 13'h00c0;
               12'b000000100010: data1 <= -13'h011c;
               12'b000000100011: data1 <= -13'h00c8;
               12'b000000100100: data1 <= 13'h015b;
               12'b000000100101: data1 <= -13'h0007;
               12'b000000100110: data1 <= 13'h01d9;
               12'b000000100111: data1 <= -13'h00d2;
               12'b000000101000: data1 <= -13'h00ae;
               12'b000000101001: data1 <= 13'h05f2;
               12'b000000101010: data1 <= 13'h004f;
               12'b000000101011: data1 <= 13'h0047;
               12'b000000101100: data1 <= 13'h00a2;
               12'b000000101101: data1 <= -13'h0025;
               12'b000000101110: data1 <= 13'h0007;
               12'b000000101111: data1 <= 13'h007b;
               12'b000000110000: data1 <= -13'h0142;
               12'b000000110001: data1 <= 13'h0008;
               12'b000000110010: data1 <= 13'h006e;
               12'b000000110011: data1 <= -13'h00b8;

endmodule: featureThreshold_rom
