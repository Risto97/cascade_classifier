module sqrt_rom
  #(
     W_DATA = 11,
     DEPTH = 64,
     W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input ena,
     input [W_ADDR-1:0] addra,
     output [W_DATA-1:0] doa

     );

     logic [W_DATA-1:0] mem [DEPTH-1:0];

     always_ff @(posedge clk)
        begin
           if(ena)
              doa = mem[addra];
        end

     initial begin
         mem[0] = 11'h00;
         mem[1] = 11'h80;
         mem[2] = 11'hb5;
         mem[3] = 11'hdd;
         mem[4] = 11'h100;
         mem[5] = 11'h11e;
         mem[6] = 11'h139;
         mem[7] = 11'h152;
         mem[8] = 11'h16a;
         mem[9] = 11'h180;
         mem[10] = 11'h194;
         mem[11] = 11'h1a8;
         mem[12] = 11'h1bb;
         mem[13] = 11'h1cd;
         mem[14] = 11'h1de;
         mem[15] = 11'h1ef;
         mem[16] = 11'h200;
         mem[17] = 11'h20f;
         mem[18] = 11'h21f;
         mem[19] = 11'h22d;
         mem[20] = 11'h23c;
         mem[21] = 11'h24a;
         mem[22] = 11'h258;
         mem[23] = 11'h265;
         mem[24] = 11'h273;
         mem[25] = 11'h280;
         mem[26] = 11'h28c;
         mem[27] = 11'h299;
         mem[28] = 11'h2a5;
         mem[29] = 11'h2b1;
         mem[30] = 11'h2bd;
         mem[31] = 11'h2c8;
         mem[32] = 11'h2d4;
         mem[33] = 11'h2df;
         mem[34] = 11'h2ea;
         mem[35] = 11'h2f5;
         mem[36] = 11'h300;
         mem[37] = 11'h30a;
         mem[38] = 11'h315;
         mem[39] = 11'h31f;
         mem[40] = 11'h329;
         mem[41] = 11'h333;
         mem[42] = 11'h33d;
         mem[43] = 11'h347;
         mem[44] = 11'h351;
         mem[45] = 11'h35a;
         mem[46] = 11'h364;
         mem[47] = 11'h36d;
         mem[48] = 11'h376;
         mem[49] = 11'h380;
         mem[50] = 11'h389;
         mem[51] = 11'h392;
         mem[52] = 11'h39b;
         mem[53] = 11'h3a3;
         mem[54] = 11'h3ac;
         mem[55] = 11'h3b5;
         mem[56] = 11'h3bd;
         mem[57] = 11'h3c6;
         mem[58] = 11'h3ce;
         mem[59] = 11'h3d7;
         mem[60] = 11'h3df;
         mem[61] = 11'h3e7;
         mem[62] = 11'h3ef;
         mem[63] = 11'h3f7;
         mem[64] = 11'h400;
         mem[65] = 11'h407;
         mem[66] = 11'h40f;
         mem[67] = 11'h417;
         mem[68] = 11'h41f;
         mem[69] = 11'h427;
         mem[70] = 11'h42e;
         mem[71] = 11'h436;
         mem[72] = 11'h43e;
         mem[73] = 11'h445;
         mem[74] = 11'h44d;
         mem[75] = 11'h454;
         mem[76] = 11'h45b;
         mem[77] = 11'h463;
         mem[78] = 11'h46a;
         mem[79] = 11'h471;
         mem[80] = 11'h478;
         mem[81] = 11'h480;
         mem[82] = 11'h487;
         mem[83] = 11'h48e;
         mem[84] = 11'h495;
         mem[85] = 11'h49c;
         mem[86] = 11'h4a3;
         mem[87] = 11'h4a9;
         mem[88] = 11'h4b0;
         mem[89] = 11'h4b7;
         mem[90] = 11'h4be;
         mem[91] = 11'h4c5;
         mem[92] = 11'h4cb;
         mem[93] = 11'h4d2;
         mem[94] = 11'h4d9;
         mem[95] = 11'h4df;
         mem[96] = 11'h4e6;
         mem[97] = 11'h4ec;
         mem[98] = 11'h4f3;
         mem[99] = 11'h4f9;
         mem[100] = 11'h500;
         mem[101] = 11'h506;
         mem[102] = 11'h50c;
         mem[103] = 11'h513;
         mem[104] = 11'h519;
         mem[105] = 11'h51f;
         mem[106] = 11'h525;
         mem[107] = 11'h52c;
         mem[108] = 11'h532;
         mem[109] = 11'h538;
         mem[110] = 11'h53e;
         mem[111] = 11'h544;
         mem[112] = 11'h54a;
         mem[113] = 11'h550;
         mem[114] = 11'h556;
         mem[115] = 11'h55c;
         mem[116] = 11'h562;
         mem[117] = 11'h568;
         mem[118] = 11'h56e;
         mem[119] = 11'h574;
         mem[120] = 11'h57a;
         mem[121] = 11'h580;
         mem[122] = 11'h585;
         mem[123] = 11'h58b;
         mem[124] = 11'h591;
         mem[125] = 11'h597;
         mem[126] = 11'h59c;
         mem[127] = 11'h5a2;
         mem[128] = 11'h5a8;
         mem[129] = 11'h5ad;
         mem[130] = 11'h5b3;
         mem[131] = 11'h5b9;
         mem[132] = 11'h5be;
         mem[133] = 11'h5c4;
         mem[134] = 11'h5c9;
         mem[135] = 11'h5cf;
         mem[136] = 11'h5d4;
         mem[137] = 11'h5da;
         mem[138] = 11'h5df;
         mem[139] = 11'h5e5;
         mem[140] = 11'h5ea;
         mem[141] = 11'h5ef;
         mem[142] = 11'h5f5;
         mem[143] = 11'h5fa;
         mem[144] = 11'h600;
         mem[145] = 11'h605;
         mem[146] = 11'h60a;
         mem[147] = 11'h60f;
         mem[148] = 11'h615;
         mem[149] = 11'h61a;
         mem[150] = 11'h61f;
         mem[151] = 11'h624;
         mem[152] = 11'h62a;
         mem[153] = 11'h62f;
         mem[154] = 11'h634;
         mem[155] = 11'h639;
         mem[156] = 11'h63e;
         mem[157] = 11'h643;
         mem[158] = 11'h648;
         mem[159] = 11'h64e;
         mem[160] = 11'h653;
         mem[161] = 11'h658;
         mem[162] = 11'h65d;
         mem[163] = 11'h662;
         mem[164] = 11'h667;
         mem[165] = 11'h66c;
         mem[166] = 11'h671;
         mem[167] = 11'h676;
         mem[168] = 11'h67b;
         mem[169] = 11'h680;
         mem[170] = 11'h684;
         mem[171] = 11'h689;
         mem[172] = 11'h68e;
         mem[173] = 11'h693;
         mem[174] = 11'h698;
         mem[175] = 11'h69d;
         mem[176] = 11'h6a2;
         mem[177] = 11'h6a6;
         mem[178] = 11'h6ab;
         mem[179] = 11'h6b0;
         mem[180] = 11'h6b5;
         mem[181] = 11'h6ba;
         mem[182] = 11'h6be;
         mem[183] = 11'h6c3;
         mem[184] = 11'h6c8;
         mem[185] = 11'h6cc;
         mem[186] = 11'h6d1;
         mem[187] = 11'h6d6;
         mem[188] = 11'h6db;
         mem[189] = 11'h6df;
         mem[190] = 11'h6e4;
         mem[191] = 11'h6e8;
         mem[192] = 11'h6ed;
         mem[193] = 11'h6f2;
         mem[194] = 11'h6f6;
         mem[195] = 11'h6fb;
         mem[196] = 11'h700;
         mem[197] = 11'h704;
         mem[198] = 11'h709;
         mem[199] = 11'h70d;
         mem[200] = 11'h712;
         mem[201] = 11'h716;
         mem[202] = 11'h71b;
         mem[203] = 11'h71f;
         mem[204] = 11'h724;
         mem[205] = 11'h728;
         mem[206] = 11'h72d;
         mem[207] = 11'h731;
         mem[208] = 11'h736;
         mem[209] = 11'h73a;
         mem[210] = 11'h73e;
         mem[211] = 11'h743;
         mem[212] = 11'h747;
         mem[213] = 11'h74c;
         mem[214] = 11'h750;
         mem[215] = 11'h754;
         mem[216] = 11'h759;
         mem[217] = 11'h75d;
         mem[218] = 11'h761;
         mem[219] = 11'h766;
         mem[220] = 11'h76a;
         mem[221] = 11'h76e;
         mem[222] = 11'h773;
         mem[223] = 11'h777;
         mem[224] = 11'h77b;
         mem[225] = 11'h780;
         mem[226] = 11'h784;
         mem[227] = 11'h788;
         mem[228] = 11'h78c;
         mem[229] = 11'h790;
         mem[230] = 11'h795;
         mem[231] = 11'h799;
         mem[232] = 11'h79d;
         mem[233] = 11'h7a1;
         mem[234] = 11'h7a6;
         mem[235] = 11'h7aa;
         mem[236] = 11'h7ae;
         mem[237] = 11'h7b2;
         mem[238] = 11'h7b6;
         mem[239] = 11'h7ba;
         mem[240] = 11'h7be;
         mem[241] = 11'h7c3;
         mem[242] = 11'h7c7;
         mem[243] = 11'h7cb;
         mem[244] = 11'h7cf;
         mem[245] = 11'h7d3;
         mem[246] = 11'h7d7;
         mem[247] = 11'h7db;
         mem[248] = 11'h7df;
         mem[249] = 11'h7e3;
         mem[250] = 11'h7e7;
         mem[251] = 11'h7eb;
         mem[252] = 11'h7ef;
         mem[253] = 11'h7f3;
         mem[254] = 11'h7f7;
         mem[255] = 11'h7fb;
     end


endmodule: sqrt_rom
