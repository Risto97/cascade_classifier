module sqrt_rom
  #(
     parameter W_DATA = 16,
     parameter W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1

     );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               8'b00000000: data1 <= 16'h0000;
               8'b00000001: data1 <= 16'h0b50;
               8'b00000010: data1 <= 16'h1000;
               8'b00000011: data1 <= 16'h1398;
               8'b00000100: data1 <= 16'h16a0;
               8'b00000101: data1 <= 16'h194c;
               8'b00000110: data1 <= 16'h1bb6;
               8'b00000111: data1 <= 16'h1dee;
               8'b00001000: data1 <= 16'h2000;
               8'b00001001: data1 <= 16'h21f0;
               8'b00001010: data1 <= 16'h23c6;
               8'b00001011: data1 <= 16'h2585;
               8'b00001100: data1 <= 16'h2731;
               8'b00001101: data1 <= 16'h28ca;
               8'b00001110: data1 <= 16'h2a54;
               8'b00001111: data1 <= 16'h2bd1;
               8'b00010000: data1 <= 16'h2d41;
               8'b00010001: data1 <= 16'h2ea5;
               8'b00010010: data1 <= 16'h3000;
               8'b00010011: data1 <= 16'h3150;
               8'b00010100: data1 <= 16'h3298;
               8'b00010101: data1 <= 16'h33d8;
               8'b00010110: data1 <= 16'h3510;
               8'b00010111: data1 <= 16'h3642;
               8'b00011000: data1 <= 16'h376c;
               8'b00011001: data1 <= 16'h3891;
               8'b00011010: data1 <= 16'h39b0;
               8'b00011011: data1 <= 16'h3ac9;
               8'b00011100: data1 <= 16'h3bdd;
               8'b00011101: data1 <= 16'h3ced;
               8'b00011110: data1 <= 16'h3df7;
               8'b00011111: data1 <= 16'h3efd;
               8'b00100000: data1 <= 16'h4000;
               8'b00100001: data1 <= 16'h40fe;
               8'b00100010: data1 <= 16'h41f8;
               8'b00100011: data1 <= 16'h42ee;
               8'b00100100: data1 <= 16'h43e1;
               8'b00100101: data1 <= 16'h44d1;
               8'b00100110: data1 <= 16'h45be;
               8'b00100111: data1 <= 16'h46a7;
               8'b00101000: data1 <= 16'h478d;
               8'b00101001: data1 <= 16'h4871;
               8'b00101010: data1 <= 16'h4952;
               8'b00101011: data1 <= 16'h4a30;
               8'b00101100: data1 <= 16'h4b0b;
               8'b00101101: data1 <= 16'h4be5;
               8'b00101110: data1 <= 16'h4cbb;
               8'b00101111: data1 <= 16'h4d90;
               8'b00110000: data1 <= 16'h4e62;
               8'b00110001: data1 <= 16'h4f32;
               8'b00110010: data1 <= 16'h5000;
               8'b00110011: data1 <= 16'h50cb;
               8'b00110100: data1 <= 16'h5195;
               8'b00110101: data1 <= 16'h525d;
               8'b00110110: data1 <= 16'h5323;
               8'b00110111: data1 <= 16'h53e7;
               8'b00111000: data1 <= 16'h54a9;
               8'b00111001: data1 <= 16'h556a;
               8'b00111010: data1 <= 16'h5629;
               8'b00111011: data1 <= 16'h56e6;
               8'b00111100: data1 <= 16'h57a2;
               8'b00111101: data1 <= 16'h585c;
               8'b00111110: data1 <= 16'h5915;
               8'b00111111: data1 <= 16'h59cc;
               8'b01000000: data1 <= 16'h5a82;
               8'b01000001: data1 <= 16'h5b36;
               8'b01000010: data1 <= 16'h5be9;
               8'b01000011: data1 <= 16'h5c9b;
               8'b01000100: data1 <= 16'h5d4b;
               8'b01000101: data1 <= 16'h5dfa;
               8'b01000110: data1 <= 16'h5ea8;
               8'b01000111: data1 <= 16'h5f54;
               8'b01001000: data1 <= 16'h6000;
               8'b01001001: data1 <= 16'h60aa;
               8'b01001010: data1 <= 16'h6152;
               8'b01001011: data1 <= 16'h61fa;
               8'b01001100: data1 <= 16'h62a1;
               8'b01001101: data1 <= 16'h6347;
               8'b01001110: data1 <= 16'h63eb;
               8'b01001111: data1 <= 16'h648e;
               8'b01010000: data1 <= 16'h6531;
               8'b01010001: data1 <= 16'h65d2;
               8'b01010010: data1 <= 16'h6673;
               8'b01010011: data1 <= 16'h6712;
               8'b01010100: data1 <= 16'h67b1;
               8'b01010101: data1 <= 16'h684e;
               8'b01010110: data1 <= 16'h68eb;
               8'b01010111: data1 <= 16'h6986;
               8'b01011000: data1 <= 16'h6a21;
               8'b01011001: data1 <= 16'h6abb;
               8'b01011010: data1 <= 16'h6b54;
               8'b01011011: data1 <= 16'h6bed;
               8'b01011100: data1 <= 16'h6c84;
               8'b01011101: data1 <= 16'h6d1a;
               8'b01011110: data1 <= 16'h6db0;
               8'b01011111: data1 <= 16'h6e45;
               8'b01100000: data1 <= 16'h6ed9;
               8'b01100001: data1 <= 16'h6f6d;
               8'b01100010: data1 <= 16'h7000;
               8'b01100011: data1 <= 16'h7091;
               8'b01100100: data1 <= 16'h7123;
               8'b01100101: data1 <= 16'h71b3;
               8'b01100110: data1 <= 16'h7243;
               8'b01100111: data1 <= 16'h72d2;
               8'b01101000: data1 <= 16'h7360;
               8'b01101001: data1 <= 16'h73ee;
               8'b01101010: data1 <= 16'h747b;
               8'b01101011: data1 <= 16'h7507;
               8'b01101100: data1 <= 16'h7593;
               8'b01101101: data1 <= 16'h761e;
               8'b01101110: data1 <= 16'h76a8;
               8'b01101111: data1 <= 16'h7732;
               8'b01110000: data1 <= 16'h77bb;
               8'b01110001: data1 <= 16'h7844;
               8'b01110010: data1 <= 16'h78cc;
               8'b01110011: data1 <= 16'h7953;
               8'b01110100: data1 <= 16'h79da;
               8'b01110101: data1 <= 16'h7a60;
               8'b01110110: data1 <= 16'h7ae5;
               8'b01110111: data1 <= 16'h7b6b;
               8'b01111000: data1 <= 16'h7bef;
               8'b01111001: data1 <= 16'h7c73;
               8'b01111010: data1 <= 16'h7cf6;
               8'b01111011: data1 <= 16'h7d79;
               8'b01111100: data1 <= 16'h7dfb;
               8'b01111101: data1 <= 16'h7e7d;
               8'b01111110: data1 <= 16'h7efe;
               8'b01111111: data1 <= 16'h7f7f;
               8'b10000000: data1 <= 16'h8000;
               8'b10000001: data1 <= 16'h807f;
               8'b10000010: data1 <= 16'h80ff;
               8'b10000011: data1 <= 16'h817d;
               8'b10000100: data1 <= 16'h81fc;
               8'b10000101: data1 <= 16'h8279;
               8'b10000110: data1 <= 16'h82f7;
               8'b10000111: data1 <= 16'h8374;
               8'b10001000: data1 <= 16'h83f0;
               8'b10001001: data1 <= 16'h846c;
               8'b10001010: data1 <= 16'h84e7;
               8'b10001011: data1 <= 16'h8562;
               8'b10001100: data1 <= 16'h85dd;
               8'b10001101: data1 <= 16'h8657;
               8'b10001110: data1 <= 16'h86d1;
               8'b10001111: data1 <= 16'h874a;
               8'b10010000: data1 <= 16'h87c3;
               8'b10010001: data1 <= 16'h883c;
               8'b10010010: data1 <= 16'h88b4;
               8'b10010011: data1 <= 16'h892b;
               8'b10010100: data1 <= 16'h89a3;
               8'b10010101: data1 <= 16'h8a19;
               8'b10010110: data1 <= 16'h8a90;
               8'b10010111: data1 <= 16'h8b06;
               8'b10011000: data1 <= 16'h8b7c;
               8'b10011001: data1 <= 16'h8bf1;
               8'b10011010: data1 <= 16'h8c66;
               8'b10011011: data1 <= 16'h8cda;
               8'b10011100: data1 <= 16'h8d4e;
               8'b10011101: data1 <= 16'h8dc2;
               8'b10011110: data1 <= 16'h8e36;
               8'b10011111: data1 <= 16'h8ea9;
               8'b10100000: data1 <= 16'h8f1b;
               8'b10100001: data1 <= 16'h8f8e;
               8'b10100010: data1 <= 16'h9000;
               8'b10100011: data1 <= 16'h9071;
               8'b10100100: data1 <= 16'h90e2;
               8'b10100101: data1 <= 16'h9153;
               8'b10100110: data1 <= 16'h91c4;
               8'b10100111: data1 <= 16'h9234;
               8'b10101000: data1 <= 16'h92a4;
               8'b10101001: data1 <= 16'h9314;
               8'b10101010: data1 <= 16'h9383;
               8'b10101011: data1 <= 16'h93f2;
               8'b10101100: data1 <= 16'h9460;
               8'b10101101: data1 <= 16'h94cf;
               8'b10101110: data1 <= 16'h953c;
               8'b10101111: data1 <= 16'h95aa;
               8'b10110000: data1 <= 16'h9617;
               8'b10110001: data1 <= 16'h9684;
               8'b10110010: data1 <= 16'h96f1;
               8'b10110011: data1 <= 16'h975d;
               8'b10110100: data1 <= 16'h97ca;
               8'b10110101: data1 <= 16'h9835;
               8'b10110110: data1 <= 16'h98a1;
               8'b10110111: data1 <= 16'h990c;
               8'b10111000: data1 <= 16'h9977;
               8'b10111001: data1 <= 16'h99e2;
               8'b10111010: data1 <= 16'h9a4c;
               8'b10111011: data1 <= 16'h9ab6;
               8'b10111100: data1 <= 16'h9b20;
               8'b10111101: data1 <= 16'h9b89;
               8'b10111110: data1 <= 16'h9bf2;
               8'b10111111: data1 <= 16'h9c5b;
               8'b11000000: data1 <= 16'h9cc4;
               8'b11000001: data1 <= 16'h9d2c;
               8'b11000010: data1 <= 16'h9d94;
               8'b11000011: data1 <= 16'h9dfc;
               8'b11000100: data1 <= 16'h9e64;
               8'b11000101: data1 <= 16'h9ecb;
               8'b11000110: data1 <= 16'h9f32;
               8'b11000111: data1 <= 16'h9f99;
               8'b11001000: data1 <= 16'ha000;
               8'b11001001: data1 <= 16'ha066;
               8'b11001010: data1 <= 16'ha0cc;
               8'b11001011: data1 <= 16'ha132;
               8'b11001100: data1 <= 16'ha197;
               8'b11001101: data1 <= 16'ha1fc;
               8'b11001110: data1 <= 16'ha261;
               8'b11001111: data1 <= 16'ha2c6;
               8'b11010000: data1 <= 16'ha32b;
               8'b11010001: data1 <= 16'ha38f;
               8'b11010010: data1 <= 16'ha3f3;
               8'b11010011: data1 <= 16'ha457;
               8'b11010100: data1 <= 16'ha4ba;
               8'b11010101: data1 <= 16'ha51e;
               8'b11010110: data1 <= 16'ha581;
               8'b11010111: data1 <= 16'ha5e4;
               8'b11011000: data1 <= 16'ha646;
               8'b11011001: data1 <= 16'ha6a9;
               8'b11011010: data1 <= 16'ha70b;
               8'b11011011: data1 <= 16'ha76d;
               8'b11011100: data1 <= 16'ha7cf;
               8'b11011101: data1 <= 16'ha830;
               8'b11011110: data1 <= 16'ha892;
               8'b11011111: data1 <= 16'ha8f3;
               8'b11100000: data1 <= 16'ha953;
               8'b11100001: data1 <= 16'ha9b4;
               8'b11100010: data1 <= 16'haa15;
               8'b11100011: data1 <= 16'haa75;
               8'b11100100: data1 <= 16'haad5;
               8'b11100101: data1 <= 16'hab35;
               8'b11100110: data1 <= 16'hab94;
               8'b11100111: data1 <= 16'habf4;
               8'b11101000: data1 <= 16'hac53;
               8'b11101001: data1 <= 16'hacb2;
               8'b11101010: data1 <= 16'had11;
               8'b11101011: data1 <= 16'had6f;
               8'b11101100: data1 <= 16'hadcd;
               8'b11101101: data1 <= 16'hae2c;
               8'b11101110: data1 <= 16'hae8a;
               8'b11101111: data1 <= 16'haee7;
               8'b11110000: data1 <= 16'haf45;
               8'b11110001: data1 <= 16'hafa2;
               8'b11110010: data1 <= 16'hb000;
               8'b11110011: data1 <= 16'hb05c;
               8'b11110100: data1 <= 16'hb0b9;
               8'b11110101: data1 <= 16'hb116;
               8'b11110110: data1 <= 16'hb172;
               8'b11110111: data1 <= 16'hb1cf;
               8'b11111000: data1 <= 16'hb22b;
               8'b11111001: data1 <= 16'hb286;
               8'b11111010: data1 <= 16'hb2e2;
               8'b11111011: data1 <= 16'hb33e;
               8'b11111100: data1 <= 16'hb399;
               8'b11111101: data1 <= 16'hb3f4;
               8'b11111110: data1 <= 16'hb44f;
               8'b11111111: data1 <= 16'hb4aa;
               default: data1 <= 0;
           endcase
        end

endmodule: sqrt_rom
