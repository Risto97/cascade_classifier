module rect1_rom
  #(
     parameter W_DATA = 20,
     parameter W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );
     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               12'b000000000000: data1 <=  20'h2d583;
               12'b000000000001: data1 <=  20'h1b887;
               12'b000000000010: data1 <=  20'h4be43;
               12'b000000000011: data1 <=  20'h7f122;
               12'b000000000100: data1 <=  20'h20853;
               12'b000000000101: data1 <=  20'h52d88;
               12'b000000000110: data1 <=  20'h46183;
               12'b000000000111: data1 <=  20'h79885;
               12'b000000001000: data1 <=  20'h13ce3;
               12'b000000001001: data1 <=  20'h33982;
               12'b000000001010: data1 <=  20'h1b887;
               12'b000000001011: data1 <=  20'h4b664;
               12'b000000001100: data1 <=  20'h0e903;
               12'b000000001101: data1 <=  20'h59cc5;
               12'b000000001110: data1 <=  20'h461c5;
               12'b000000001111: data1 <=  20'h141c3;
               12'b000000010000: data1 <=  20'h48c66;
               12'b000000010001: data1 <=  20'h2184a;
               12'b000000010010: data1 <=  20'h3504a;
               12'b000000010011: data1 <=  20'h20449;
               12'b000000010100: data1 <=  20'h0504b;
               12'b000000010101: data1 <=  20'h2790d;
               12'b000000010110: data1 <=  20'h28449;
               12'b000000010111: data1 <=  20'h7ed42;
               12'b000000011000: data1 <=  20'h529c6;
               12'b000000011001: data1 <=  20'h14d03;
               12'b000000011010: data1 <=  20'h461e3;
               12'b000000011011: data1 <=  20'h538a7;
               12'b000000011100: data1 <=  20'h2204a;
               12'b000000011101: data1 <=  20'h4c866;
               12'b000000011110: data1 <=  20'h858c3;
               12'b000000011111: data1 <=  20'h335a2;
               12'b000000100000: data1 <=  20'h0ac6f;
               12'b000000100001: data1 <=  20'h0746f;
               12'b000000100010: data1 <=  20'h3410f;
               12'b000000100011: data1 <=  20'h26ce6;
               12'b000000100100: data1 <=  20'h64aa4;
               12'b000000100101: data1 <=  20'h08c4a;
               12'b000000100110: data1 <=  20'h51d4a;
               12'b000000100111: data1 <=  20'h06c4d;
               12'b000000101000: data1 <=  20'h1184d;
               12'b000000101001: data1 <=  20'h22173;
               12'b000000101010: data1 <=  20'h1e049;
               12'b000000101011: data1 <=  20'h1344b;
               12'b000000101100: data1 <=  20'h09449;
               12'b000000101101: data1 <=  20'h2be61;
               12'b000000101110: data1 <=  20'h09449;
               12'b000000101111: data1 <=  20'h08c49;
               12'b000000110000: data1 <=  20'h224e7;
               12'b000000110001: data1 <=  20'h45241;
               12'b000000110010: data1 <=  20'h5584b;
               12'b000000110011: data1 <=  20'h2bcc3;
               12'b000000110100: data1 <=  20'h2d583;
               12'b000000110101: data1 <=  20'h21c86;
               12'b000000110110: data1 <=  20'h08505;
               12'b000000110111: data1 <=  20'h4c242;
               12'b000000111000: data1 <=  20'h6acc3;
               12'b000000111001: data1 <=  20'h1784d;
               12'b000000111010: data1 <=  20'h1384d;
               12'b000000111011: data1 <=  20'h08517;
               12'b000000111100: data1 <=  20'h45104;
               12'b000000111101: data1 <=  20'h5b067;
               12'b000000111110: data1 <=  20'h4bd03;
               12'b000000111111: data1 <=  20'h33982;
               12'b000001000000: data1 <=  20'h534c6;
               12'b000001000001: data1 <=  20'h6e122;
               12'b000001000010: data1 <=  20'h70e41;
               12'b000001000011: data1 <=  20'h3fa06;
               12'b000001000100: data1 <=  20'h06c54;
               12'b000001000101: data1 <=  20'h07241;
               12'b000001000110: data1 <=  20'h1f947;
               12'b000001000111: data1 <=  20'h4c5c4;
               12'b000001001000: data1 <=  20'h6b0e3;
               12'b000001001001: data1 <=  20'h6dd22;
               12'b000001001010: data1 <=  20'h6a922;
               12'b000001001011: data1 <=  20'h29485;
               12'b000001001100: data1 <=  20'h208e7;
               12'b000001001101: data1 <=  20'h02885;
               12'b000001001110: data1 <=  20'h150c3;
               12'b000001001111: data1 <=  20'h28449;
               12'b000001010000: data1 <=  20'h02449;
               12'b000001010001: data1 <=  20'h28849;
               12'b000001010010: data1 <=  20'h28049;
               12'b000001010011: data1 <=  20'h344c4;
               12'b000001010100: data1 <=  20'h14583;
               12'b000001010101: data1 <=  20'h02106;
               12'b000001010110: data1 <=  20'h45e04;
               12'b000001010111: data1 <=  20'h28466;
               12'b000001011000: data1 <=  20'h7f103;
               12'b000001011001: data1 <=  20'h28449;
               12'b000001011010: data1 <=  20'h538a4;
               12'b000001011011: data1 <=  20'h28449;
               12'b000001011100: data1 <=  20'h28449;
               12'b000001011101: data1 <=  20'h72cc6;
               12'b000001011110: data1 <=  20'h90241;
               12'b000001011111: data1 <=  20'h4d885;
               12'b000001100000: data1 <=  20'h4c905;
               12'b000001100001: data1 <=  20'h33d42;
               12'b000001100010: data1 <=  20'h64142;
               12'b000001100011: data1 <=  20'h78641;
               12'b000001100100: data1 <=  20'h0cec1;
               12'b000001100101: data1 <=  20'h6be41;
               12'b000001100110: data1 <=  20'h1a46f;
               12'b000001100111: data1 <=  20'h1e04a;
               12'b000001101000: data1 <=  20'h1984a;
               12'b000001101001: data1 <=  20'h67143;
               12'b000001101010: data1 <=  20'h4c089;
               12'b000001101011: data1 <=  20'h03849;
               12'b000001101100: data1 <=  20'h40866;
               12'b000001101101: data1 <=  20'h364c3;
               12'b000001101110: data1 <=  20'h320c3;
               12'b000001101111: data1 <=  20'h03849;
               12'b000001110000: data1 <=  20'h02049;
               12'b000001110001: data1 <=  20'h66122;
               12'b000001110010: data1 <=  20'h70922;
               12'b000001110011: data1 <=  20'h3504a;
               12'b000001110100: data1 <=  20'h790c3;
               12'b000001110101: data1 <=  20'h45681;
               12'b000001110110: data1 <=  20'h38d26;
               12'b000001110111: data1 <=  20'h00d38;
               12'b000001111000: data1 <=  20'h26ce5;
               12'b000001111001: data1 <=  20'h22ca6;
               12'b000001111010: data1 <=  20'h204c6;
               12'b000001111011: data1 <=  20'h5ee41;
               12'b000001111100: data1 <=  20'h6bd04;
               12'b000001111101: data1 <=  20'h77a43;
               12'b000001111110: data1 <=  20'h00c66;
               12'b000001111111: data1 <=  20'h28092;
               12'b000010000000: data1 <=  20'h0844e;
               12'b000010000001: data1 <=  20'h13a61;
               12'b000010000010: data1 <=  20'h3516d;
               12'b000010000011: data1 <=  20'h46d62;
               12'b000010000100: data1 <=  20'h4c4aa;
               12'b000010000101: data1 <=  20'h68086;
               12'b000010000110: data1 <=  20'h65086;
               12'b000010000111: data1 <=  20'h240a4;
               12'b000010001000: data1 <=  20'h0e904;
               12'b000010001001: data1 <=  20'h40182;
               12'b000010001010: data1 <=  20'h21c66;
               12'b000010001011: data1 <=  20'h7f4c3;
               12'b000010001100: data1 <=  20'h4b2c5;
               12'b000010001101: data1 <=  20'h1a223;
               12'b000010001110: data1 <=  20'h2184a;
               12'b000010001111: data1 <=  20'h0ac68;
               12'b000010010000: data1 <=  20'h07067;
               12'b000010010001: data1 <=  20'h04876;
               12'b000010010010: data1 <=  20'h00c76;
               12'b000010010011: data1 <=  20'h2fc90;
               12'b000010010100: data1 <=  20'h4ba62;
               12'b000010010101: data1 <=  20'h538c4;
               12'b000010010110: data1 <=  20'h6ae22;
               12'b000010010111: data1 <=  20'h5b067;
               12'b000010011000: data1 <=  20'h26c85;
               12'b000010011001: data1 <=  20'h3686b;
               12'b000010011010: data1 <=  20'h32c6b;
               12'b000010011011: data1 <=  20'h5fd49;
               12'b000010011100: data1 <=  20'h59467;
               12'b000010011101: data1 <=  20'h59908;
               12'b000010011110: data1 <=  20'h4112e;
               12'b000010011111: data1 <=  20'h614c3;
               12'b000010100000: data1 <=  20'h01ca8;
               12'b000010100001: data1 <=  20'h03466;
               12'b000010100010: data1 <=  20'h15d04;
               12'b000010100011: data1 <=  20'h03466;
               12'b000010100100: data1 <=  20'h06942;
               12'b000010100101: data1 <=  20'h03466;
               12'b000010100110: data1 <=  20'h02066;
               12'b000010100111: data1 <=  20'h7f142;
               12'b000010101000: data1 <=  20'h14c49;
               12'b000010101001: data1 <=  20'h21182;
               12'b000010101010: data1 <=  20'h44e41;
               12'b000010101011: data1 <=  20'h452c1;
               12'b000010101100: data1 <=  20'h47088;
               12'b000010101101: data1 <=  20'h47c66;
               12'b000010101110: data1 <=  20'h47066;
               12'b000010101111: data1 <=  20'h4cd62;
               12'b000010110000: data1 <=  20'h51582;
               12'b000010110001: data1 <=  20'h1c566;
               12'b000010110010: data1 <=  20'h03151;
               12'b000010110011: data1 <=  20'h03838;
               12'b000010110100: data1 <=  20'h02438;
               12'b000010110101: data1 <=  20'h09c36;
               12'b000010110110: data1 <=  20'h08836;
               12'b000010110111: data1 <=  20'h2a032;
               12'b000010111000: data1 <=  20'h65922;
               12'b000010111001: data1 <=  20'h67522;
               12'b000010111010: data1 <=  20'h77a41;
               12'b000010111011: data1 <=  20'h1c489;
               12'b000010111100: data1 <=  20'h70a41;
               12'b000010111101: data1 <=  20'h0e0c4;
               12'b000010111110: data1 <=  20'h465c3;
               12'b000010111111: data1 <=  20'h21c66;
               12'b000011000000: data1 <=  20'h53cc8;
               12'b000011000001: data1 <=  20'h1a070;
               12'b000011000010: data1 <=  20'h14243;
               12'b000011000011: data1 <=  20'h790a4;
               12'b000011000100: data1 <=  20'h05049;
               12'b000011000101: data1 <=  20'h06e41;
               12'b000011000110: data1 <=  20'h91261;
               12'b000011000111: data1 <=  20'h00849;
               12'b000011001000: data1 <=  20'h4c666;
               12'b000011001001: data1 <=  20'h06c49;
               12'b000011001010: data1 <=  20'h228e6;
               12'b000011001011: data1 <=  20'h0ca81;
               12'b000011001100: data1 <=  20'h132c1;
               12'b000011001101: data1 <=  20'h454e3;
               12'b000011001110: data1 <=  20'h4e562;
               12'b000011001111: data1 <=  20'h4b162;
               12'b000011010000: data1 <=  20'h2e84b;
               12'b000011010001: data1 <=  20'h08c66;
               12'b000011010010: data1 <=  20'h2e885;
               12'b000011010011: data1 <=  20'h40186;
               12'b000011010100: data1 <=  20'h2a0c5;
               12'b000011010101: data1 <=  20'h64e41;
               12'b000011010110: data1 <=  20'h368c3;
               12'b000011010111: data1 <=  20'h1f903;
               12'b000011011000: data1 <=  20'h03449;
               12'b000011011001: data1 <=  20'h19187;
               12'b000011011010: data1 <=  20'h0344d;
               12'b000011011011: data1 <=  20'h0244d;
               12'b000011011100: data1 <=  20'h28c49;
               12'b000011011101: data1 <=  20'h2e449;
               12'b000011011110: data1 <=  20'h7a122;
               12'b000011011111: data1 <=  20'h710e3;
               12'b000011100000: data1 <=  20'h73922;
               12'b000011100001: data1 <=  20'h7e4a4;
               12'b000011100010: data1 <=  20'h614a9;
               12'b000011100011: data1 <=  20'h26a02;
               12'b000011100100: data1 <=  20'h33d42;
               12'b000011100101: data1 <=  20'h58caa;
               12'b000011100110: data1 <=  20'h3b4a7;
               12'b000011100111: data1 <=  20'h27c49;
               12'b000011101000: data1 <=  20'h2ca41;
               12'b000011101001: data1 <=  20'h44e41;
               12'b000011101010: data1 <=  20'h67122;
               12'b000011101011: data1 <=  20'h268e3;
               12'b000011101100: data1 <=  20'h03432;
               12'b000011101101: data1 <=  20'h02832;
               12'b000011101110: data1 <=  20'h2e4aa;
               12'b000011101111: data1 <=  20'h7f0e4;
               12'b000011110000: data1 <=  20'h5a0a9;
               12'b000011110001: data1 <=  20'h0c983;
               12'b000011110010: data1 <=  20'h09564;
               12'b000011110011: data1 <=  20'h13de3;
               12'b000011110100: data1 <=  20'h02113;
               12'b000011110101: data1 <=  20'h86123;
               12'b000011110110: data1 <=  20'h2e0a4;
               12'b000011110111: data1 <=  20'h2e4a4;
               12'b000011111000: data1 <=  20'h37068;
               12'b000011111001: data1 <=  20'h5e142;
               12'b000011111010: data1 <=  20'h6dd42;
               12'b000011111011: data1 <=  20'h13a03;
               12'b000011111100: data1 <=  20'h488e5;
               12'b000011111101: data1 <=  20'h0904d;
               12'b000011111110: data1 <=  20'h10c6e;
               12'b000011111111: data1 <=  20'h584c5;
               12'b000100000000: data1 <=  20'h33d42;
               12'b000100000001: data1 <=  20'h0d86e;
               12'b000100000010: data1 <=  20'h348a4;
               12'b000100000011: data1 <=  20'h6c505;
               12'b000100000100: data1 <=  20'h488a4;
               12'b000100000101: data1 <=  20'h07066;
               12'b000100000110: data1 <=  20'h670c3;
               12'b000100000111: data1 <=  20'h658c3;
               12'b000100001000: data1 <=  20'h5b068;
               12'b000100001001: data1 <=  20'h57da2;
               12'b000100001010: data1 <=  20'h09849;
               12'b000100001011: data1 <=  20'h02866;
               12'b000100001100: data1 <=  20'h0f869;
               12'b000100001101: data1 <=  20'h0ec69;
               12'b000100001110: data1 <=  20'h7e982;
               12'b000100001111: data1 <=  20'h27c49;
               12'b000100010000: data1 <=  20'h2d8c3;
               12'b000100010001: data1 <=  20'h40907;
               12'b000100010010: data1 <=  20'h33d44;
               12'b000100010011: data1 <=  20'h190c3;
               12'b000100010100: data1 <=  20'h10434;
               12'b000100010101: data1 <=  20'h258c3;
               12'b000100010110: data1 <=  20'h16835;
               12'b000100010111: data1 <=  20'h02037;
               12'b000100011000: data1 <=  20'h42522;
               12'b000100011001: data1 <=  20'h3e922;
               12'b000100011010: data1 <=  20'h66122;
               12'b000100011011: data1 <=  20'h64122;
               12'b000100011100: data1 <=  20'h40cc4;
               12'b000100011101: data1 <=  20'h02113;
               12'b000100011110: data1 <=  20'h2e106;
               12'b000100011111: data1 <=  20'h2884a;
               12'b000100100000: data1 <=  20'h3b4a6;
               12'b000100100001: data1 <=  20'h01833;
               12'b000100100010: data1 <=  20'h0404a;
               12'b000100100011: data1 <=  20'h00866;
               12'b000100100100: data1 <=  20'h4b301;
               12'b000100100101: data1 <=  20'h45da2;
               12'b000100100110: data1 <=  20'h470c3;
               12'b000100100111: data1 <=  20'h57a02;
               12'b000100101000: data1 <=  20'h624c3;
               12'b000100101001: data1 <=  20'h5dcc3;
               12'b000100101010: data1 <=  20'h2dca4;
               12'b000100101011: data1 <=  20'h2e449;
               12'b000100101100: data1 <=  20'h03449;
               12'b000100101101: data1 <=  20'h02449;
               12'b000100101110: data1 <=  20'h1644f;
               12'b000100101111: data1 <=  20'h14c4f;
               12'b000100110000: data1 <=  20'h1cd22;
               12'b000100110001: data1 <=  20'h40867;
               12'b000100110010: data1 <=  20'h790c5;
               12'b000100110011: data1 <=  20'h6c0a4;
               12'b000100110100: data1 <=  20'h54c68;
               12'b000100110101: data1 <=  20'h71241;
               12'b000100110110: data1 <=  20'h78261;
               12'b000100110111: data1 <=  20'h02c49;
               12'b000100111000: data1 <=  20'h1c432;
               12'b000100111001: data1 <=  20'h1b832;
               12'b000100111010: data1 <=  20'h150c9;
               12'b000100111011: data1 <=  20'h0844e;
               12'b000100111100: data1 <=  20'h79d23;
               12'b000100111101: data1 <=  20'h13148;
               12'b000100111110: data1 <=  20'h23066;
               12'b000100111111: data1 <=  20'h0cd68;
               12'b000101000000: data1 <=  20'h794a5;
               12'b000101000001: data1 <=  20'h8a641;
               12'b000101000010: data1 <=  20'h5a84a;
               12'b000101000011: data1 <=  20'h0e904;
               12'b000101000100: data1 <=  20'h2d583;
               12'b000101000101: data1 <=  20'h28085;
               12'b000101000110: data1 <=  20'h4c5c4;
               12'b000101000111: data1 <=  20'h58885;
               12'b000101001000: data1 <=  20'h540a7;
               12'b000101001001: data1 <=  20'h59468;
               12'b000101001010: data1 <=  20'h2e0c8;
               12'b000101001011: data1 <=  20'h19a81;
               12'b000101001100: data1 <=  20'h58662;
               12'b000101001101: data1 <=  20'h28049;
               12'b000101001110: data1 <=  20'h2986e;
               12'b000101001111: data1 <=  20'h3a84c;
               12'b000101010000: data1 <=  20'h2ac69;
               12'b000101010001: data1 <=  20'h25869;
               12'b000101010010: data1 <=  20'h23cc3;
               12'b000101010011: data1 <=  20'h7dde2;
               12'b000101010100: data1 <=  20'h23cc3;
               12'b000101010101: data1 <=  20'h1f4c3;
               12'b000101010110: data1 <=  20'h46241;
               12'b000101010111: data1 <=  20'h0e182;
               12'b000101011000: data1 <=  20'h03049;
               12'b000101011001: data1 <=  20'h02849;
               12'b000101011010: data1 <=  20'h5b522;
               12'b000101011011: data1 <=  20'h32da2;
               12'b000101011100: data1 <=  20'h5b522;
               12'b000101011101: data1 <=  20'h2086f;
               12'b000101011110: data1 <=  20'h34c66;
               12'b000101011111: data1 <=  20'h53467;
               12'b000101100000: data1 <=  20'h5b522;
               12'b000101100001: data1 <=  20'h4d4a4;
               12'b000101100010: data1 <=  20'h09853;
               12'b000101100011: data1 <=  20'h08853;
               12'b000101100100: data1 <=  20'h4f8c3;
               12'b000101100101: data1 <=  20'h89e41;
               12'b000101100110: data1 <=  20'h67943;
               12'b000101100111: data1 <=  20'h51962;
               12'b000101101000: data1 <=  20'h28903;
               12'b000101101001: data1 <=  20'h0052b;
               12'b000101101010: data1 <=  20'h2f487;
               12'b000101101011: data1 <=  20'h1906a;
               12'b000101101100: data1 <=  20'h04449;
               12'b000101101101: data1 <=  20'h01449;
               12'b000101101110: data1 <=  20'h4f866;
               12'b000101101111: data1 <=  20'h4bc66;
               12'b000101110000: data1 <=  20'h5b522;
               12'b000101110001: data1 <=  20'h57922;
               12'b000101110010: data1 <=  20'h5ee61;
               12'b000101110011: data1 <=  20'h58261;
               12'b000101110100: data1 <=  20'h6dd42;
               12'b000101110101: data1 <=  20'h018a6;
               12'b000101110110: data1 <=  20'h0b466;
               12'b000101110111: data1 <=  20'h06866;
               12'b000101111000: data1 <=  20'h6e4c3;
               12'b000101111001: data1 <=  20'h3a126;
               12'b000101111010: data1 <=  20'h2ec86;
               12'b000101111011: data1 <=  20'h1a1c4;
               12'b000101111100: data1 <=  20'h28849;
               12'b000101111101: data1 <=  20'h408c3;
               12'b000101111110: data1 <=  20'h6e122;
               12'b000101111111: data1 <=  20'h080f7;
               12'b000110000000: data1 <=  20'h46622;
               12'b000110000001: data1 <=  20'h25d66;
               12'b000110000010: data1 <=  20'h6bda2;
               12'b000110000011: data1 <=  20'h6a522;
               12'b000110000100: data1 <=  20'h2f0a4;
               12'b000110000101: data1 <=  20'h600c3;
               12'b000110000110: data1 <=  20'h350c3;
               12'b000110000111: data1 <=  20'h59904;
               12'b000110001000: data1 <=  20'h68066;
               12'b000110001001: data1 <=  20'h19301;
               12'b000110001010: data1 <=  20'h7a542;
               12'b000110001011: data1 <=  20'h530c3;
               12'b000110001100: data1 <=  20'h14243;
               12'b000110001101: data1 <=  20'h26a03;
               12'b000110001110: data1 <=  20'h48c66;
               12'b000110001111: data1 <=  20'h2d4c4;
               12'b000110010000: data1 <=  20'h28849;
               12'b000110010001: data1 <=  20'h34c4a;
               12'b000110010010: data1 <=  20'h60849;
               12'b000110010011: data1 <=  20'h09535;
               12'b000110010100: data1 <=  20'h338c7;
               12'b000110010101: data1 <=  20'h21c49;
               12'b000110010110: data1 <=  20'h0e904;
               12'b000110010111: data1 <=  20'h484a4;
               12'b000110011000: data1 <=  20'h460a4;
               12'b000110011001: data1 <=  20'h28449;
               12'b000110011010: data1 <=  20'h07071;
               12'b000110011011: data1 <=  20'h19e63;
               12'b000110011100: data1 <=  20'h714c3;
               12'b000110011101: data1 <=  20'h1e053;
               12'b000110011110: data1 <=  20'h654a7;
               12'b000110011111: data1 <=  20'h2f0a6;
               12'b000110100000: data1 <=  20'h2d4a6;
               12'b000110100001: data1 <=  20'h0f866;
               12'b000110100010: data1 <=  20'h7f0e4;
               12'b000110100011: data1 <=  20'h59d22;
               12'b000110100100: data1 <=  20'h0f066;
               12'b000110100101: data1 <=  20'h0344e;
               12'b000110100110: data1 <=  20'h0244e;
               12'b000110100111: data1 <=  20'h6dd22;
               12'b000110101000: data1 <=  20'h340c5;
               12'b000110101001: data1 <=  20'h17c4b;
               12'b000110101010: data1 <=  20'h4c967;
               12'b000110101011: data1 <=  20'h304c3;
               12'b000110101100: data1 <=  20'h33d22;
               12'b000110101101: data1 <=  20'h304c3;
               12'b000110101110: data1 <=  20'h2bcc3;
               12'b000110101111: data1 <=  20'h27d22;
               12'b000110110000: data1 <=  20'h8fe61;
               12'b000110110001: data1 <=  20'h6e8c3;
               12'b000110110010: data1 <=  20'h6a8c3;
               12'b000110110011: data1 <=  20'h48449;
               12'b000110110100: data1 <=  20'h46c49;
               12'b000110110101: data1 <=  20'h3a8c7;
               12'b000110110110: data1 <=  20'h6c8c5;
               12'b000110110111: data1 <=  20'h03849;
               12'b000110111000: data1 <=  20'h02049;
               12'b000110111001: data1 <=  20'h72241;
               12'b000110111010: data1 <=  20'h70e41;
               12'b000110111011: data1 <=  20'h4d966;
               12'b000110111100: data1 <=  20'h26ce3;
               12'b000110111101: data1 <=  20'h26de2;
               12'b000110111110: data1 <=  20'h066c1;
               12'b000110111111: data1 <=  20'h02118;
               12'b000111000000: data1 <=  20'h60524;
               12'b000111000001: data1 <=  20'h46583;
               12'b000111000010: data1 <=  20'h650e4;
               12'b000111000011: data1 <=  20'h0f963;
               12'b000111000100: data1 <=  20'h800e3;
               12'b000111000101: data1 <=  20'h03188;
               12'b000111000110: data1 <=  20'h52122;
               12'b000111000111: data1 <=  20'h456c1;
               12'b000111001000: data1 <=  20'h2d564;
               12'b000111001001: data1 <=  20'h358c3;
               12'b000111001010: data1 <=  20'h38702;
               12'b000111001011: data1 <=  20'h04ca5;
               12'b000111001100: data1 <=  20'h000a5;
               12'b000111001101: data1 <=  20'h09582;
               12'b000111001110: data1 <=  20'h70a41;
               12'b000111001111: data1 <=  20'h61103;
               12'b000111010000: data1 <=  20'h5e903;
               12'b000111010001: data1 <=  20'h6be41;
               12'b000111010010: data1 <=  20'h70aa5;
               12'b000111010011: data1 <=  20'h03c58;
               12'b000111010100: data1 <=  20'h1b44b;
               12'b000111010101: data1 <=  20'h22466;
               12'b000111010110: data1 <=  20'h57c4a;
               12'b000111010111: data1 <=  20'h03c58;
               12'b000111011000: data1 <=  20'h01c58;
               12'b000111011001: data1 <=  20'h30867;
               12'b000111011010: data1 <=  20'h2d44c;
               12'b000111011011: data1 <=  20'h2150e;
               12'b000111011100: data1 <=  20'h5f142;
               12'b000111011101: data1 <=  20'h03849;
               12'b000111011110: data1 <=  20'h2c467;
               12'b000111011111: data1 <=  20'h1106f;
               12'b000111100000: data1 <=  20'h0d049;
               12'b000111100001: data1 <=  20'h10ca7;
               12'b000111100010: data1 <=  20'h28832;
               12'b000111100011: data1 <=  20'h22ca6;
               12'b000111100100: data1 <=  20'h2804a;
               12'b000111100101: data1 <=  20'h03849;
               12'b000111100110: data1 <=  20'h14467;
               12'b000111100111: data1 <=  20'h2d4e3;
               12'b000111101000: data1 <=  20'h2e886;
               12'b000111101001: data1 <=  20'h544e6;
               12'b000111101010: data1 <=  20'h28049;
               12'b000111101011: data1 <=  20'h6e4c3;
               12'b000111101100: data1 <=  20'h0184d;
               12'b000111101101: data1 <=  20'h0ece3;
               12'b000111101110: data1 <=  20'h334a4;
               12'b000111101111: data1 <=  20'h34885;
               12'b000111110000: data1 <=  20'h340a4;
               12'b000111110001: data1 <=  20'h14563;
               12'b000111110010: data1 <=  20'h28085;
               12'b000111110011: data1 <=  20'h02105;
               12'b000111110100: data1 <=  20'h4b6e2;
               12'b000111110101: data1 <=  20'h858c3;
               12'b000111110110: data1 <=  20'h32ea2;
               12'b000111110111: data1 <=  20'h1fc4c;
               12'b000111111000: data1 <=  20'h2e485;
               12'b000111111001: data1 <=  20'h4d105;
               12'b000111111010: data1 <=  20'h2e4ac;
               12'b000111111011: data1 <=  20'h76d42;
               12'b000111111100: data1 <=  20'h80922;
               12'b000111111101: data1 <=  20'h59cc8;
               12'b000111111110: data1 <=  20'h80922;
               12'b000111111111: data1 <=  20'h7d522;
               12'b001000000000: data1 <=  20'h48922;
               12'b001000000001: data1 <=  20'h44d22;
               12'b001000000010: data1 <=  20'h17849;
               12'b001000000011: data1 <=  20'h71241;
               12'b001000000100: data1 <=  20'h6b2a2;
               12'b001000000101: data1 <=  20'h7f4c3;
               12'b001000000110: data1 <=  20'h2a0c3;
               12'b001000000111: data1 <=  20'h258c3;
               12'b001000001000: data1 <=  20'h03105;
               12'b001000001001: data1 <=  20'h008a8;
               12'b001000001010: data1 <=  20'h038a5;
               12'b001000001011: data1 <=  20'h014a5;
               12'b001000001100: data1 <=  20'h1746a;
               12'b001000001101: data1 <=  20'h460c3;
               12'b001000001110: data1 <=  20'h05832;
               12'b001000001111: data1 <=  20'h02049;
               12'b001000010000: data1 <=  20'h34c67;
               12'b001000010001: data1 <=  20'h4cc85;
               12'b001000010010: data1 <=  20'h05832;
               12'b001000010011: data1 <=  20'h28849;
               12'b001000010100: data1 <=  20'h10522;
               12'b001000010101: data1 <=  20'h12f01;
               12'b001000010110: data1 <=  20'h2f049;
               12'b001000010111: data1 <=  20'h27c4a;
               12'b001000011000: data1 <=  20'h09c4c;
               12'b001000011001: data1 <=  20'h40186;
               12'b001000011010: data1 <=  20'h16435;
               12'b001000011011: data1 <=  20'h20d84;
               12'b001000011100: data1 <=  20'h19e44;
               12'b001000011101: data1 <=  20'h07241;
               12'b001000011110: data1 <=  20'h54582;
               12'b001000011111: data1 <=  20'h22449;
               12'b001000100000: data1 <=  20'h09849;
               12'b001000100001: data1 <=  20'h0e856;
               12'b001000100010: data1 <=  20'h43887;
               12'b001000100011: data1 <=  20'h39205;
               12'b001000100100: data1 <=  20'h43887;
               12'b001000100101: data1 <=  20'h3e887;
               12'b001000100110: data1 <=  20'h6cd63;
               12'b001000100111: data1 <=  20'h2dd09;
               12'b001000101000: data1 <=  20'h09850;
               12'b001000101001: data1 <=  20'h08850;
               12'b001000101010: data1 <=  20'h22904;
               12'b001000101011: data1 <=  20'h4b0c3;
               12'b001000101100: data1 <=  20'h6be41;
               12'b001000101101: data1 <=  20'h5e8c3;
               12'b001000101110: data1 <=  20'h66122;
               12'b001000101111: data1 <=  20'h51c85;
               12'b001000110000: data1 <=  20'h48866;
               12'b001000110001: data1 <=  20'h26641;
               12'b001000110010: data1 <=  20'h2404b;
               12'b001000110011: data1 <=  20'h2004b;
               12'b001000110100: data1 <=  20'h0b049;
               12'b001000110101: data1 <=  20'h07049;
               12'b001000110110: data1 <=  20'h5ed29;
               12'b001000110111: data1 <=  20'h46582;
               12'b001000111000: data1 <=  20'h1cd22;
               12'b001000111001: data1 <=  20'h19122;
               12'b001000111010: data1 <=  20'h04451;
               12'b001000111011: data1 <=  20'h01451;
               12'b001000111100: data1 <=  20'h78d22;
               12'b001000111101: data1 <=  20'h46466;
               12'b001000111110: data1 <=  20'h335c6;
               12'b001000111111: data1 <=  20'h34866;
               12'b001001000000: data1 <=  20'h4d9c5;
               12'b001001000001: data1 <=  20'h4b1c5;
               12'b001001000010: data1 <=  20'h10522;
               12'b001001000011: data1 <=  20'h0c922;
               12'b001001000100: data1 <=  20'h2904e;
               12'b001001000101: data1 <=  20'h2e849;
               12'b001001000110: data1 <=  20'h2904f;
               12'b001001000111: data1 <=  20'h2784f;
               12'b001001001000: data1 <=  20'h16889;
               12'b001001001001: data1 <=  20'h00c75;
               12'b001001001010: data1 <=  20'h54104;
               12'b001001001011: data1 <=  20'h2d4a6;
               12'b001001001100: data1 <=  20'h28849;
               12'b001001001101: data1 <=  20'h12cc3;
               12'b001001001110: data1 <=  20'h5ea41;
               12'b001001001111: data1 <=  20'h58485;
               12'b001001010000: data1 <=  20'h4e182;
               12'b001001010001: data1 <=  20'h0cc34;
               12'b001001010010: data1 <=  20'h684a4;
               12'b001001010011: data1 <=  20'h648a4;
               12'b001001010100: data1 <=  20'h14943;
               12'b001001010101: data1 <=  20'h02103;
               12'b001001010110: data1 <=  20'h3f5e2;
               12'b001001010111: data1 <=  20'h21c86;
               12'b001001011000: data1 <=  20'h655c3;
               12'b001001011001: data1 <=  20'h79885;
               12'b001001011010: data1 <=  20'h26467;
               12'b001001011011: data1 <=  20'h04866;
               12'b001001011100: data1 <=  20'h0d641;
               12'b001001011101: data1 <=  20'h4d5c6;
               12'b001001011110: data1 <=  20'h00c66;
               12'b001001011111: data1 <=  20'h48066;
               12'b001001100000: data1 <=  20'h7f103;
               12'b001001100001: data1 <=  20'h48067;
               12'b001001100010: data1 <=  20'h58942;
               12'b001001100011: data1 <=  20'h48066;
               12'b001001100100: data1 <=  20'h46c67;
               12'b001001100101: data1 <=  20'h33d64;
               12'b001001100110: data1 <=  20'h6bd42;
               12'b001001100111: data1 <=  20'h04049;
               12'b001001101000: data1 <=  20'h01849;
               12'b001001101001: data1 <=  20'h2e885;
               12'b001001101010: data1 <=  20'h06681;
               12'b001001101011: data1 <=  20'h80542;
               12'b001001101100: data1 <=  20'h2d06b;
               12'b001001101101: data1 <=  20'h6cd43;
               12'b001001101110: data1 <=  20'h0f049;
               12'b001001101111: data1 <=  20'h164a4;
               12'b001001110000: data1 <=  20'h270c3;
               12'b001001110001: data1 <=  20'h35085;
               12'b001001110010: data1 <=  20'h4cc88;
               12'b001001110011: data1 <=  20'h40922;
               12'b001001110100: data1 <=  20'h209c3;
               12'b001001110101: data1 <=  20'h7de64;
               12'b001001110110: data1 <=  20'h014a8;
               12'b001001110111: data1 <=  20'h0dd12;
               12'b001001111000: data1 <=  20'h46d0b;
               12'b001001111001: data1 <=  20'h13925;
               12'b001001111010: data1 <=  20'h6aa41;
               12'b001001111011: data1 <=  20'h71e41;
               12'b001001111100: data1 <=  20'h5e122;
               12'b001001111101: data1 <=  20'h57ee5;
               12'b001001111110: data1 <=  20'h32e41;
               12'b001001111111: data1 <=  20'h338c3;
               12'b001010000000: data1 <=  20'h0e436;
               12'b001010000001: data1 <=  20'h7a542;
               12'b001010000010: data1 <=  20'h7d542;
               12'b001010000011: data1 <=  20'h1604c;
               12'b001010000100: data1 <=  20'h28849;
               12'b001010000101: data1 <=  20'h03449;
               12'b001010000110: data1 <=  20'h02449;
               12'b001010000111: data1 <=  20'h42466;
               12'b001010001000: data1 <=  20'h46069;
               12'b001010001001: data1 <=  20'h23033;
               12'b001010001010: data1 <=  20'h33922;
               12'b001010001011: data1 <=  20'h23033;
               12'b001010001100: data1 <=  20'h258c3;
               12'b001010001101: data1 <=  20'h8ae41;
               12'b001010001110: data1 <=  20'h404c4;
               12'b001010001111: data1 <=  20'h1d485;
               12'b001010010000: data1 <=  20'h34866;
               12'b001010010001: data1 <=  20'h3c068;
               12'b001010010010: data1 <=  20'h3e8a4;
               12'b001010010011: data1 <=  20'h290e3;
               12'b001010010100: data1 <=  20'h21433;
               12'b001010010101: data1 <=  20'h1c4b4;
               12'b001010010110: data1 <=  20'h1a8b4;
               12'b001010010111: data1 <=  20'h41c66;
               12'b001010011000: data1 <=  20'h40866;
               12'b001010011001: data1 <=  20'h10c67;
               12'b001010011010: data1 <=  20'h0d867;
               12'b001010011011: data1 <=  20'h1c067;
               12'b001010011100: data1 <=  20'h1bc49;
               12'b001010011101: data1 <=  20'h1bc8a;
               12'b001010011110: data1 <=  20'h1b48a;
               12'b001010011111: data1 <=  20'h7f142;
               12'b001010100000: data1 <=  20'h7d6a2;
               12'b001010100001: data1 <=  20'h0ecc6;
               12'b001010100010: data1 <=  20'h0ecc6;
               12'b001010100011: data1 <=  20'h23cc3;
               12'b001010100100: data1 <=  20'h46cc3;
               12'b001010100101: data1 <=  20'h38e82;
               12'b001010100110: data1 <=  20'h1f4c3;
               12'b001010100111: data1 <=  20'h5c085;
               12'b001010101000: data1 <=  20'h58085;
               12'b001010101001: data1 <=  20'h4554d;
               12'b001010101010: data1 <=  20'h3b4c5;
               12'b001010101011: data1 <=  20'h28d03;
               12'b001010101100: data1 <=  20'h83922;
               12'b001010101101: data1 <=  20'h22085;
               12'b001010101110: data1 <=  20'h200e6;
               12'b001010101111: data1 <=  20'h1c066;
               12'b001010110000: data1 <=  20'h2c661;
               12'b001010110001: data1 <=  20'h55cc3;
               12'b001010110010: data1 <=  20'h32e41;
               12'b001010110011: data1 <=  20'h12049;
               12'b001010110100: data1 <=  20'h77681;
               12'b001010110101: data1 <=  20'h3eec1;
               12'b001010110110: data1 <=  20'h0c849;
               12'b001010110111: data1 <=  20'h04c57;
               12'b001010111000: data1 <=  20'h13873;
               12'b001010111001: data1 <=  20'h11849;
               12'b001010111010: data1 <=  20'h2bd42;
               12'b001010111011: data1 <=  20'h034c6;
               12'b001010111100: data1 <=  20'h12d83;
               12'b001010111101: data1 <=  20'h79485;
               12'b001010111110: data1 <=  20'h59885;
               12'b001010111111: data1 <=  20'h58a23;
               12'b001011000000: data1 <=  20'h1fd24;
               12'b001011000001: data1 <=  20'h290e3;
               12'b001011000010: data1 <=  20'h264e3;
               12'b001011000011: data1 <=  20'h23832;
               12'b001011000100: data1 <=  20'h20c32;
               12'b001011000101: data1 <=  20'h4d9c2;
               12'b001011000110: data1 <=  20'h4c122;
               12'b001011000111: data1 <=  20'h13643;
               12'b001011001000: data1 <=  20'h15488;
               12'b001011001001: data1 <=  20'h07885;
               12'b001011001010: data1 <=  20'h47ce4;
               12'b001011001011: data1 <=  20'h57ac2;
               12'b001011001100: data1 <=  20'h48885;
               12'b001011001101: data1 <=  20'h460e4;
               12'b001011001110: data1 <=  20'h7f122;
               12'b001011001111: data1 <=  20'h196c2;
               12'b001011010000: data1 <=  20'h17851;
               12'b001011010001: data1 <=  20'h46d09;
               12'b001011010010: data1 <=  20'h05066;
               12'b001011010011: data1 <=  20'h02449;
               12'b001011010100: data1 <=  20'h48926;
               12'b001011010101: data1 <=  20'h90641;
               12'b001011010110: data1 <=  20'h428c3;
               12'b001011010111: data1 <=  20'h06c4b;
               12'b001011011000: data1 <=  20'h0504a;
               12'b001011011001: data1 <=  20'h13851;
               12'b001011011010: data1 <=  20'h6e122;
               12'b001011011011: data1 <=  20'h64103;
               12'b001011011100: data1 <=  20'h4f0c4;
               12'b001011011101: data1 <=  20'h4b8c4;
               12'b001011011110: data1 <=  20'h2e485;
               12'b001011011111: data1 <=  20'h25e61;
               12'b001011100000: data1 <=  20'h35867;
               12'b001011100001: data1 <=  20'h45983;
               12'b001011100010: data1 <=  20'h2ca41;
               12'b001011100011: data1 <=  20'h28086;
               12'b001011100100: data1 <=  20'h3912e;
               12'b001011100101: data1 <=  20'h00849;
               12'b001011100110: data1 <=  20'h22452;
               12'b001011100111: data1 <=  20'h21c52;
               12'b001011101000: data1 <=  20'h2244a;
               12'b001011101001: data1 <=  20'h1bc4b;
               12'b001011101010: data1 <=  20'h6b641;
               12'b001011101011: data1 <=  20'h6a681;
               12'b001011101100: data1 <=  20'h538c4;
               12'b001011101101: data1 <=  20'h6c504;
               12'b001011101110: data1 <=  20'h67466;
               12'b001011101111: data1 <=  20'h398e7;
               12'b001011110000: data1 <=  20'h03185;
               12'b001011110001: data1 <=  20'h4b641;
               12'b001011110010: data1 <=  20'h3d0a4;
               12'b001011110011: data1 <=  20'h384a4;
               12'b001011110100: data1 <=  20'h2a889;
               12'b001011110101: data1 <=  20'h25889;
               12'b001011110110: data1 <=  20'h23cc6;
               12'b001011110111: data1 <=  20'h27c49;
               12'b001011111000: data1 <=  20'h5404b;
               12'b001011111001: data1 <=  20'h1f4c6;
               12'b001011111010: data1 <=  20'h132e1;
               12'b001011111011: data1 <=  20'h64661;
               12'b001011111100: data1 <=  20'h7a162;
               12'b001011111101: data1 <=  20'h52485;
               12'b001011111110: data1 <=  20'h418a4;
               12'b001011111111: data1 <=  20'h39523;
               12'b001100000000: data1 <=  20'h67d22;
               12'b001100000001: data1 <=  20'h57d22;
               12'b001100000010: data1 <=  20'h41d44;
               12'b001100000011: data1 <=  20'h01472;
               12'b001100000100: data1 <=  20'h48c6a;
               12'b001100000101: data1 <=  20'h0dc85;
               12'b001100000110: data1 <=  20'h1b8e6;
               12'b001100000111: data1 <=  20'h01ca7;
               12'b001100001000: data1 <=  20'h79d82;
               12'b001100001001: data1 <=  20'h322e2;
               12'b001100001010: data1 <=  20'h42c85;
               12'b001100001011: data1 <=  20'h6a641;
               12'b001100001100: data1 <=  20'h74522;
               12'b001100001101: data1 <=  20'h70922;
               12'b001100001110: data1 <=  20'h48066;
               12'b001100001111: data1 <=  20'h46c66;
               12'b001100010000: data1 <=  20'h15d83;
               12'b001100010001: data1 <=  20'h1fe41;
               12'b001100010010: data1 <=  20'h03182;
               12'b001100010011: data1 <=  20'h6aa41;
               12'b001100010100: data1 <=  20'h6e122;
               12'b001100010101: data1 <=  20'h6a522;
               12'b001100010110: data1 <=  20'h72241;
               12'b001100010111: data1 <=  20'h3484a;
               12'b001100011000: data1 <=  20'h28849;
               12'b001100011001: data1 <=  20'h4d0a4;
               12'b001100011010: data1 <=  20'h4e0c4;
               12'b001100011011: data1 <=  20'h2144b;
               12'b001100011100: data1 <=  20'h3b903;
               12'b001100011101: data1 <=  20'h38aa2;
               12'b001100011110: data1 <=  20'h48866;
               12'b001100011111: data1 <=  20'h52d64;
               12'b001100100000: data1 <=  20'h368a4;
               12'b001100100001: data1 <=  20'h34cc3;
               12'b001100100010: data1 <=  20'h47cc4;
               12'b001100100011: data1 <=  20'h44ecb;
               12'b001100100100: data1 <=  20'h284c4;
               12'b001100100101: data1 <=  20'h02c49;
               12'b001100100110: data1 <=  20'h03049;
               12'b001100100111: data1 <=  20'h14c67;
               12'b001100101000: data1 <=  20'h40cc8;
               12'b001100101001: data1 <=  20'h2e467;
               12'b001100101010: data1 <=  20'h5260a;
               12'b001100101011: data1 <=  20'h1bc4a;
               12'b001100101100: data1 <=  20'h0de02;
               12'b001100101101: data1 <=  20'h214c4;
               12'b001100101110: data1 <=  20'h03c49;
               12'b001100101111: data1 <=  20'h1c085;
               12'b001100110000: data1 <=  20'h418a4;
               12'b001100110001: data1 <=  20'h404a4;
               12'b001100110010: data1 <=  20'h47885;
               12'b001100110011: data1 <=  20'h3f485;
               12'b001100110100: data1 <=  20'h4e868;
               12'b001100110101: data1 <=  20'h85503;
               12'b001100110110: data1 <=  20'h7f4c4;
               12'b001100110111: data1 <=  20'h6a922;
               12'b001100111000: data1 <=  20'h79942;
               12'b001100111001: data1 <=  20'h72c86;
               12'b001100111010: data1 <=  20'h28866;
               12'b001100111011: data1 <=  20'h644c3;
               12'b001100111100: data1 <=  20'h72182;
               12'b001100111101: data1 <=  20'h25e81;
               12'b001100111110: data1 <=  20'h1b123;
               12'b001100111111: data1 <=  20'h83d22;
               12'b001101000000: data1 <=  20'h2e886;
               12'b001101000001: data1 <=  20'h0e486;
               12'b001101000010: data1 <=  20'h42068;
               12'b001101000011: data1 <=  20'h47085;
               12'b001101000100: data1 <=  20'h3bc66;
               12'b001101000101: data1 <=  20'h40449;
               12'b001101000110: data1 <=  20'h45ca4;
               12'b001101000111: data1 <=  20'h024e6;
               12'b001101001000: data1 <=  20'h33d42;
               12'b001101001001: data1 <=  20'h02c4f;
               12'b001101001010: data1 <=  20'h13641;
               12'b001101001011: data1 <=  20'h7f103;
               12'b001101001100: data1 <=  20'h07241;
               12'b001101001101: data1 <=  20'h02c66;
               12'b001101001110: data1 <=  20'h70a41;
               12'b001101001111: data1 <=  20'h2e485;
               12'b001101010000: data1 <=  20'h13449;
               12'b001101010001: data1 <=  20'h11849;
               12'b001101010010: data1 <=  20'h0d049;
               12'b001101010011: data1 <=  20'h09582;
               12'b001101010100: data1 <=  20'h70922;
               12'b001101010101: data1 <=  20'h61522;
               12'b001101010110: data1 <=  20'h64261;
               12'b001101010111: data1 <=  20'h22566;
               12'b001101011000: data1 <=  20'h53466;
               12'b001101011001: data1 <=  20'h13e81;
               12'b001101011010: data1 <=  20'h5a04a;
               12'b001101011011: data1 <=  20'h4e903;
               12'b001101011100: data1 <=  20'h64903;
               12'b001101011101: data1 <=  20'h35867;
               12'b001101011110: data1 <=  20'h4b903;
               12'b001101011111: data1 <=  20'h7e604;
               12'b001101100000: data1 <=  20'h2e086;
               12'b001101100001: data1 <=  20'h0f885;
               12'b001101100010: data1 <=  20'h270c3;
               12'b001101100011: data1 <=  20'h2ec49;
               12'b001101100100: data1 <=  20'h00086;
               12'b001101100101: data1 <=  20'h494c3;
               12'b001101100110: data1 <=  20'h4c466;
               12'b001101100111: data1 <=  20'h85ce3;
               12'b001101101000: data1 <=  20'h13603;
               12'b001101101001: data1 <=  20'h3b8e3;
               12'b001101101010: data1 <=  20'h46487;
               12'b001101101011: data1 <=  20'h2e849;
               12'b001101101100: data1 <=  20'h33c67;
               12'b001101101101: data1 <=  20'h68888;
               12'b001101101110: data1 <=  20'h5a44a;
               12'b001101101111: data1 <=  20'h47485;
               12'b001101110000: data1 <=  20'h516e1;
               12'b001101110001: data1 <=  20'h03c4c;
               12'b001101110010: data1 <=  20'h3f885;
               12'b001101110011: data1 <=  20'h1c542;
               12'b001101110100: data1 <=  20'h01c4c;
               12'b001101110101: data1 <=  20'h29066;
               12'b001101110110: data1 <=  20'h27466;
               12'b001101110111: data1 <=  20'h47ccd;
               12'b001101111000: data1 <=  20'h464cd;
               12'b001101111001: data1 <=  20'h68086;
               12'b001101111010: data1 <=  20'h2bea1;
               12'b001101111011: data1 <=  20'h68086;
               12'b001101111100: data1 <=  20'h58cc7;
               12'b001101111101: data1 <=  20'h46261;
               12'b001101111110: data1 <=  20'h26dc2;
               12'b001101111111: data1 <=  20'h72cc4;
               12'b001110000000: data1 <=  20'h02449;
               12'b001110000001: data1 <=  20'h22962;
               12'b001110000010: data1 <=  20'h01466;
               12'b001110000011: data1 <=  20'h0b057;
               12'b001110000100: data1 <=  20'h07057;
               12'b001110000101: data1 <=  20'h6ba41;
               12'b001110000110: data1 <=  20'h1f562;
               12'b001110000111: data1 <=  20'h6ae81;
               12'b001110001000: data1 <=  20'h209a2;
               12'b001110001001: data1 <=  20'h3896f;
               12'b001110001010: data1 <=  20'h1b8e3;
               12'b001110001011: data1 <=  20'h2dca4;
               12'b001110001100: data1 <=  20'h2e8a4;
               12'b001110001101: data1 <=  20'h1c049;
               12'b001110001110: data1 <=  20'h4c066;
               12'b001110001111: data1 <=  20'h15c85;
               12'b001110010000: data1 <=  20'h26503;
               12'b001110010001: data1 <=  20'h399c3;
               12'b001110010010: data1 <=  20'h20522;
               12'b001110010011: data1 <=  20'h1aa41;
               12'b001110010100: data1 <=  20'h28066;
               12'b001110010101: data1 <=  20'h0cb01;
               12'b001110010110: data1 <=  20'h76d42;
               12'b001110010111: data1 <=  20'h77a41;
               12'b001110011000: data1 <=  20'h1fc68;
               12'b001110011001: data1 <=  20'h33d62;
               12'b001110011010: data1 <=  20'h5298b;
               12'b001110011011: data1 <=  20'h4d885;
               12'b001110011100: data1 <=  20'h27c86;
               12'b001110011101: data1 <=  20'h494c3;
               12'b001110011110: data1 <=  20'h2e0aa;
               12'b001110011111: data1 <=  20'h22449;
               12'b001110100000: data1 <=  20'h3b04a;
               12'b001110100001: data1 <=  20'h5ac4a;
               12'b001110100010: data1 <=  20'h59c4a;
               12'b001110100011: data1 <=  20'h45e03;
               12'b001110100100: data1 <=  20'h4ba81;
               12'b001110100101: data1 <=  20'h0344d;
               12'b001110100110: data1 <=  20'h0244d;
               12'b001110100111: data1 <=  20'h088c7;
               12'b001110101000: data1 <=  20'h57cc3;
               12'b001110101001: data1 <=  20'h7f122;
               12'b001110101010: data1 <=  20'h459e2;
               12'b001110101011: data1 <=  20'h46261;
               12'b001110101100: data1 <=  20'h598e8;
               12'b001110101101: data1 <=  20'h66522;
               12'b001110101110: data1 <=  20'h44d04;
               12'b001110101111: data1 <=  20'h20e41;
               12'b001110110000: data1 <=  20'h65086;
               12'b001110110001: data1 <=  20'h61122;
               12'b001110110010: data1 <=  20'h334e7;
               12'b001110110011: data1 <=  20'h67163;
               12'b001110110100: data1 <=  20'h02c49;
               12'b001110110101: data1 <=  20'h22ca5;
               12'b001110110110: data1 <=  20'h208a5;
               12'b001110110111: data1 <=  20'h28903;
               12'b001110111000: data1 <=  20'h3e8c3;
               12'b001110111001: data1 <=  20'h43887;
               12'b001110111010: data1 <=  20'h72cc6;
               12'b001110111011: data1 <=  20'h41886;
               12'b001110111100: data1 <=  20'h02849;
               12'b001110111101: data1 <=  20'h1c888;
               12'b001110111110: data1 <=  20'h4cd42;
               12'b001110111111: data1 <=  20'h288e7;
               12'b001111000000: data1 <=  20'h4ba81;
               12'b001111000001: data1 <=  20'h68888;
               12'b001111000010: data1 <=  20'h450c5;
               12'b001111000011: data1 <=  20'h46582;
               12'b001111000100: data1 <=  20'h4e067;
               12'b001111000101: data1 <=  20'h1c888;
               12'b001111000110: data1 <=  20'h1a888;
               12'b001111000111: data1 <=  20'h3b066;
               12'b001111001000: data1 <=  20'h1f906;
               12'b001111001001: data1 <=  20'h3a868;
               12'b001111001010: data1 <=  20'h01c32;
               12'b001111001011: data1 <=  20'h684a7;
               12'b001111001100: data1 <=  20'h648a7;
               12'b001111001101: data1 <=  20'h2d943;
               12'b001111001110: data1 <=  20'h38ae6;
               12'b001111001111: data1 <=  20'h084e3;
               12'b001111010000: data1 <=  20'h28449;
               12'b001111010001: data1 <=  20'h714c3;
               12'b001111010010: data1 <=  20'h37088;
               12'b001111010011: data1 <=  20'h78d04;
               12'b001111010100: data1 <=  20'h37088;
               12'b001111010101: data1 <=  20'h32088;
               12'b001111010110: data1 <=  20'h6c505;
               12'b001111010111: data1 <=  20'h460a4;
               12'b001111011000: data1 <=  20'h0da61;
               12'b001111011001: data1 <=  20'h4d109;
               12'b001111011010: data1 <=  20'h1a9a4;
               12'b001111011011: data1 <=  20'h06701;
               12'b001111011100: data1 <=  20'h17c4b;
               12'b001111011101: data1 <=  20'h28049;
               12'b001111011110: data1 <=  20'h47cc4;
               12'b001111011111: data1 <=  20'h320c3;
               12'b001111100000: data1 <=  20'h72241;
               12'b001111100001: data1 <=  20'h64122;
               12'b001111100010: data1 <=  20'h17c49;
               12'b001111100011: data1 <=  20'h13449;
               12'b001111100100: data1 <=  20'h04873;
               12'b001111100101: data1 <=  20'h00c73;
               12'b001111100110: data1 <=  20'h48068;
               12'b001111100111: data1 <=  20'h46c68;
               12'b001111101000: data1 <=  20'h4c661;
               12'b001111101001: data1 <=  20'h7f4c4;
               12'b001111101010: data1 <=  20'h33a02;
               12'b001111101011: data1 <=  20'h02466;
               12'b001111101100: data1 <=  20'h41087;
               12'b001111101101: data1 <=  20'h451e6;
               12'b001111101110: data1 <=  20'h4dc85;
               12'b001111101111: data1 <=  20'h01c49;
               12'b001111110000: data1 <=  20'h03849;
               12'b001111110001: data1 <=  20'h208c4;
               12'b001111110010: data1 <=  20'h5ad62;
               12'b001111110011: data1 <=  20'h57aa1;
               12'b001111110100: data1 <=  20'h09486;
               12'b001111110101: data1 <=  20'h00466;
               12'b001111110110: data1 <=  20'h136a1;
               12'b001111110111: data1 <=  20'h13661;
               12'b001111111000: data1 <=  20'h43867;
               12'b001111111001: data1 <=  20'h3ec67;
               12'b001111111010: data1 <=  20'h290e7;
               12'b001111111011: data1 <=  20'h57922;
               12'b001111111100: data1 <=  20'h6e103;
               12'b001111111101: data1 <=  20'h06962;
               12'b001111111110: data1 <=  20'h53922;
               12'b001111111111: data1 <=  20'h64241;
               12'b010000000000: data1 <=  20'h6e4e3;
               12'b010000000001: data1 <=  20'h15d04;
               12'b010000000010: data1 <=  20'h274c5;
               12'b010000000011: data1 <=  20'h28449;
               12'b010000000100: data1 <=  20'h0944a;
               12'b010000000101: data1 <=  20'h08c4a;
               12'b010000000110: data1 <=  20'h744c3;
               12'b010000000111: data1 <=  20'h714c3;
               12'b010000001000: data1 <=  20'h0a433;
               12'b010000001001: data1 <=  20'h13849;
               12'b010000001010: data1 <=  20'h04033;
               12'b010000001011: data1 <=  20'h15cc4;
               12'b010000001100: data1 <=  20'h21c49;
               12'b010000001101: data1 <=  20'h01c33;
               12'b010000001110: data1 <=  20'h2e866;
               12'b010000001111: data1 <=  20'h2e8a5;
               12'b010000010000: data1 <=  20'h15c32;
               12'b010000010001: data1 <=  20'h1584c;
               12'b010000010010: data1 <=  20'h32e61;
               12'b010000010011: data1 <=  20'h32a41;
               12'b010000010100: data1 <=  20'h54522;
               12'b010000010101: data1 <=  20'h20849;
               12'b010000010110: data1 <=  20'h09d42;
               12'b010000010111: data1 <=  20'h06542;
               12'b010000011000: data1 <=  20'h60466;
               12'b010000011001: data1 <=  20'h0e908;
               12'b010000011010: data1 <=  20'h26e41;
               12'b010000011011: data1 <=  20'h60866;
               12'b010000011100: data1 <=  20'h4dc85;
               12'b010000011101: data1 <=  20'h4d485;
               12'b010000011110: data1 <=  20'h0ddc2;
               12'b010000011111: data1 <=  20'h2e485;
               12'b010000100000: data1 <=  20'h474a4;
               12'b010000100001: data1 <=  20'h3a087;
               12'b010000100010: data1 <=  20'h22563;
               12'b010000100011: data1 <=  20'h320c3;
               12'b010000100100: data1 <=  20'h79d22;
               12'b010000100101: data1 <=  20'h77661;
               12'b010000100110: data1 <=  20'h79d22;
               12'b010000100111: data1 <=  20'h70e41;
               12'b010000101000: data1 <=  20'h79d22;
               12'b010000101001: data1 <=  20'h06701;
               12'b010000101010: data1 <=  20'h0ddc2;
               12'b010000101011: data1 <=  20'h65922;
               12'b010000101100: data1 <=  20'h678c3;
               12'b010000101101: data1 <=  20'h8ada2;
               12'b010000101110: data1 <=  20'h538c4;
               12'b010000101111: data1 <=  20'h408e3;
               12'b010000110000: data1 <=  20'h34c66;
               12'b010000110001: data1 <=  20'h40067;
               12'b010000110010: data1 <=  20'h42ca4;
               12'b010000110011: data1 <=  20'h5fd03;
               12'b010000110100: data1 <=  20'h2dd22;
               12'b010000110101: data1 <=  20'h650c3;
               12'b010000110110: data1 <=  20'h79d22;
               12'b010000110111: data1 <=  20'h600c3;
               12'b010000111000: data1 <=  20'h3c4e5;
               12'b010000111001: data1 <=  20'h388e5;
               12'b010000111010: data1 <=  20'h2e871;
               12'b010000111011: data1 <=  20'h19c6a;
               12'b010000111100: data1 <=  20'h33ca4;
               12'b010000111101: data1 <=  20'h2ec49;
               12'b010000111110: data1 <=  20'h60c49;
               12'b010000111111: data1 <=  20'h32c68;
               12'b010001000000: data1 <=  20'h79d22;
               12'b010001000001: data1 <=  20'h77922;
               12'b010001000010: data1 <=  20'h09866;
               12'b010001000011: data1 <=  20'h4c485;
               12'b010001000100: data1 <=  20'h22086;
               12'b010001000101: data1 <=  20'h1b468;
               12'b010001000110: data1 <=  20'h684a4;
               12'b010001000111: data1 <=  20'h648a4;
               12'b010001001000: data1 <=  20'h03182;
               12'b010001001001: data1 <=  20'h32122;
               12'b010001001010: data1 <=  20'h1c183;
               12'b010001001011: data1 <=  20'h0dd62;
               12'b010001001100: data1 <=  20'h09562;
               12'b010001001101: data1 <=  20'h600c9;
               12'b010001001110: data1 <=  20'h45682;
               12'b010001001111: data1 <=  20'h399c7;
               12'b010001010000: data1 <=  20'h20603;
               12'b010001010001: data1 <=  20'h19a61;
               12'b010001010010: data1 <=  20'h14942;
               12'b010001010011: data1 <=  20'h57885;
               12'b010001010100: data1 <=  20'h456a1;
               12'b010001010101: data1 <=  20'h01866;
               12'b010001010110: data1 <=  20'h2d5c3;
               12'b010001010111: data1 <=  20'h09049;
               12'b010001011000: data1 <=  20'h48923;
               12'b010001011001: data1 <=  20'h2dc87;
               12'b010001011010: data1 <=  20'h90a61;
               12'b010001011011: data1 <=  20'h64a81;
               12'b010001011100: data1 <=  20'h04c4d;
               12'b010001011101: data1 <=  20'h45104;
               12'b010001011110: data1 <=  20'h6dcc3;
               12'b010001011111: data1 <=  20'h6b4c3;
               12'b010001100000: data1 <=  20'h22c4a;
               12'b010001100001: data1 <=  20'h2144a;
               12'b010001100010: data1 <=  20'h358c3;
               12'b010001100011: data1 <=  20'h330c3;
               12'b010001100100: data1 <=  20'h0e915;
               12'b010001100101: data1 <=  20'h0d44d;
               12'b010001100110: data1 <=  20'h05055;
               12'b010001100111: data1 <=  20'h19854;
               12'b010001101000: data1 <=  20'h72922;
               12'b010001101001: data1 <=  20'h02449;
               12'b010001101010: data1 <=  20'h61ce3;
               12'b010001101011: data1 <=  20'h864e3;
               12'b010001101100: data1 <=  20'h22069;
               12'b010001101101: data1 <=  20'h2244a;
               12'b010001101110: data1 <=  20'h28849;
               12'b010001101111: data1 <=  20'h21c69;
               12'b010001110000: data1 <=  20'h67942;
               12'b010001110001: data1 <=  20'h208e7;
               12'b010001110010: data1 <=  20'h368c3;
               12'b010001110011: data1 <=  20'h270c6;
               12'b010001110100: data1 <=  20'h5484a;
               12'b010001110101: data1 <=  20'h3ed44;
               12'b010001110110: data1 <=  20'h61922;
               12'b010001110111: data1 <=  20'h150c3;
               12'b010001111000: data1 <=  20'h348a7;
               12'b010001111001: data1 <=  20'h26602;
               12'b010001111010: data1 <=  20'h29903;
               12'b010001111011: data1 <=  20'h5384a;
               12'b010001111100: data1 <=  20'h61922;
               12'b010001111101: data1 <=  20'h5dd22;
               12'b010001111110: data1 <=  20'h73d22;
               12'b010001111111: data1 <=  20'h71122;
               12'b010010000000: data1 <=  20'h6ba41;
               12'b010010000001: data1 <=  20'h6aa41;
               12'b010010000010: data1 <=  20'h07a41;
               12'b010010000011: data1 <=  20'h0ce61;
               12'b010010000100: data1 <=  20'h1084b;
               12'b010010000101: data1 <=  20'h600a6;
               12'b010010000110: data1 <=  20'h1084b;
               12'b010010000111: data1 <=  20'h0e04b;
               12'b010010001000: data1 <=  20'h23cc3;
               12'b010010001001: data1 <=  20'h0cd62;
               12'b010010001010: data1 <=  20'h024ec;
               12'b010010001011: data1 <=  20'h51641;
               12'b010010001100: data1 <=  20'h10049;
               12'b010010001101: data1 <=  20'h45a41;
               12'b010010001110: data1 <=  20'h29903;
               12'b010010001111: data1 <=  20'h32e41;
               12'b010010010000: data1 <=  20'h47849;
               12'b010010010001: data1 <=  20'h34c49;
               12'b010010010010: data1 <=  20'h03c32;
               12'b010010010011: data1 <=  20'h02032;
               12'b010010010100: data1 <=  20'h29ce3;
               12'b010010010101: data1 <=  20'h7dd22;
               12'b010010010110: data1 <=  20'h77aa1;
               12'b010010010111: data1 <=  20'h258e3;
               12'b010010011000: data1 <=  20'h32ac1;
               12'b010010011001: data1 <=  20'h12d88;
               12'b010010011010: data1 <=  20'h7a122;
               12'b010010011011: data1 <=  20'h208c4;
               12'b010010011100: data1 <=  20'h288e3;
               12'b010010011101: data1 <=  20'h654e3;
               12'b010010011110: data1 <=  20'h23cc3;
               12'b010010011111: data1 <=  20'h1f4c3;
               12'b010010100000: data1 <=  20'h1c545;
               12'b010010100001: data1 <=  20'h52868;
               12'b010010100010: data1 <=  20'h088ef;
               12'b010010100011: data1 <=  20'h4e0e8;
               12'b010010100100: data1 <=  20'h2d4c4;
               12'b010010100101: data1 <=  20'h21866;
               12'b010010100110: data1 <=  20'h48066;
               12'b010010100111: data1 <=  20'h46c66;
               12'b010010101000: data1 <=  20'h20e41;
               12'b010010101001: data1 <=  20'h0d04b;
               12'b010010101010: data1 <=  20'h0504f;
               12'b010010101011: data1 <=  20'h0084d;
               12'b010010101100: data1 <=  20'h03849;
               12'b010010101101: data1 <=  20'h02049;
               12'b010010101110: data1 <=  20'h0e904;
               12'b010010101111: data1 <=  20'h54524;
               12'b010010110000: data1 <=  20'h2e0a4;
               12'b010010110001: data1 <=  20'h34cc3;
               12'b010010110010: data1 <=  20'h5ee61;
               12'b010010110011: data1 <=  20'h4108a;
               12'b010010110100: data1 <=  20'h6c522;
               12'b010010110101: data1 <=  20'h3a0a4;
               12'b010010110110: data1 <=  20'h1c087;
               12'b010010110111: data1 <=  20'h514c3;
               12'b010010111000: data1 <=  20'h368c3;
               12'b010010111001: data1 <=  20'h70903;
               12'b010010111010: data1 <=  20'h748e3;
               12'b010010111011: data1 <=  20'h7d542;
               12'b010010111100: data1 <=  20'h35143;
               12'b010010111101: data1 <=  20'h34449;
               12'b010010111110: data1 <=  20'h22488;
               12'b010010111111: data1 <=  20'h21488;
               12'b010011000000: data1 <=  20'h28849;
               12'b010011000001: data1 <=  20'h01050;
               12'b010011000010: data1 <=  20'h35cc4;
               12'b010011000011: data1 <=  20'h32cc4;
               12'b010011000100: data1 <=  20'h5b522;
               12'b010011000101: data1 <=  20'h45deb;
               12'b010011000110: data1 <=  20'h5b522;
               12'b010011000111: data1 <=  20'h57922;
               12'b010011001000: data1 <=  20'h6e122;
               12'b010011001001: data1 <=  20'h6a522;
               12'b010011001010: data1 <=  20'h03885;
               12'b010011001011: data1 <=  20'h00c50;
               12'b010011001100: data1 <=  20'h33d42;
               12'b010011001101: data1 <=  20'h6cc85;
               12'b010011001110: data1 <=  20'h27942;
               12'b010011001111: data1 <=  20'h8c922;
               12'b010011010000: data1 <=  20'h3a162;
               12'b010011010001: data1 <=  20'h000c5;
               12'b010011010010: data1 <=  20'h0a4c3;
               12'b010011010011: data1 <=  20'h72522;
               12'b010011010100: data1 <=  20'h2e4b0;
               12'b010011010101: data1 <=  20'h414cd;
               12'b010011010110: data1 <=  20'h0f8c3;
               12'b010011010111: data1 <=  20'h4bd83;
               12'b010011011000: data1 <=  20'h23503;
               12'b010011011001: data1 <=  20'h1f503;
               12'b010011011010: data1 <=  20'h12d8b;
               12'b010011011011: data1 <=  20'h51485;
               12'b010011011100: data1 <=  20'h79485;
               12'b010011011101: data1 <=  20'h3ac87;
               12'b010011011110: data1 <=  20'h2cde3;
               12'b010011011111: data1 <=  20'h08506;
               12'b010011100000: data1 <=  20'h59ca8;
               12'b010011100001: data1 <=  20'h858c3;
               12'b010011100010: data1 <=  20'h46466;
               12'b010011100011: data1 <=  20'h28449;
               12'b010011100100: data1 <=  20'h27868;
               12'b010011100101: data1 <=  20'h1a281;
               12'b010011100110: data1 <=  20'h408c3;
               12'b010011100111: data1 <=  20'h6c142;
               12'b010011101000: data1 <=  20'h19449;
               12'b010011101001: data1 <=  20'h03c49;
               12'b010011101010: data1 <=  20'h01c49;
               12'b010011101011: data1 <=  20'h03449;
               12'b010011101100: data1 <=  20'h2e066;
               12'b010011101101: data1 <=  20'h07241;
               12'b010011101110: data1 <=  20'h3e942;
               12'b010011101111: data1 <=  20'h34886;
               12'b010011110000: data1 <=  20'h20c66;
               12'b010011110001: data1 <=  20'h03d2b;
               12'b010011110010: data1 <=  20'h0012b;
               12'b010011110011: data1 <=  20'h1184b;
               12'b010011110100: data1 <=  20'h0d04b;
               12'b010011110101: data1 <=  20'h03449;
               12'b010011110110: data1 <=  20'h06681;
               12'b010011110111: data1 <=  20'h13681;
               12'b010011111000: data1 <=  20'h45241;
               12'b010011111001: data1 <=  20'h430c3;
               12'b010011111010: data1 <=  20'h12ec3;
               12'b010011111011: data1 <=  20'h29cc3;
               12'b010011111100: data1 <=  20'h3e8c3;
               12'b010011111101: data1 <=  20'h32302;
               12'b010011111110: data1 <=  20'h0d04a;
               12'b010011111111: data1 <=  20'h28849;
               12'b010100000000: data1 <=  20'h02449;
               12'b010100000001: data1 <=  20'h04449;
               12'b010100000010: data1 <=  20'h01449;
               12'b010100000011: data1 <=  20'h7a922;
               12'b010100000100: data1 <=  20'h70a41;
               12'b010100000101: data1 <=  20'h67d22;
               12'b010100000110: data1 <=  20'h6a6e2;
               12'b010100000111: data1 <=  20'h65641;
               12'b010100001000: data1 <=  20'h64122;
               12'b010100001001: data1 <=  20'h35485;
               12'b010100001010: data1 <=  20'h2dca6;
               12'b010100001011: data1 <=  20'h35485;
               12'b010100001100: data1 <=  20'h0206c;
               12'b010100001101: data1 <=  20'h35485;
               12'b010100001110: data1 <=  20'h21c49;
               12'b010100001111: data1 <=  20'h28849;
               12'b010100010000: data1 <=  20'h2e8c4;
               12'b010100010001: data1 <=  20'h35485;
               12'b010100010010: data1 <=  20'h33c85;
               12'b010100010011: data1 <=  20'h42067;
               12'b010100010100: data1 <=  20'h22473;
               12'b010100010101: data1 <=  20'h4e0c3;
               12'b010100010110: data1 <=  20'h38923;
               12'b010100010111: data1 <=  20'h5c885;
               12'b010100011000: data1 <=  20'h38564;
               12'b010100011001: data1 <=  20'h740c3;
               12'b010100011010: data1 <=  20'h25949;
               12'b010100011011: data1 <=  20'h28d46;
               12'b010100011100: data1 <=  20'h640a4;
               12'b010100011101: data1 <=  20'h6be41;
               12'b010100011110: data1 <=  20'h4b261;
               12'b010100011111: data1 <=  20'h3bcc3;
               12'b010100100000: data1 <=  20'h2c162;
               12'b010100100001: data1 <=  20'h41ce4;
               12'b010100100010: data1 <=  20'h3f963;
               12'b010100100011: data1 <=  20'h42ca4;
               12'b010100100100: data1 <=  20'h4c467;
               12'b010100100101: data1 <=  20'h6e4c3;
               12'b010100100110: data1 <=  20'h64cc4;
               12'b010100100111: data1 <=  20'h678c3;
               12'b010100101000: data1 <=  20'h02849;
               12'b010100101001: data1 <=  20'h09057;
               12'b010100101010: data1 <=  20'h70922;
               12'b010100101011: data1 <=  20'h71a41;
               12'b010100101100: data1 <=  20'h399a7;
               12'b010100101101: data1 <=  20'h04c86;
               12'b010100101110: data1 <=  20'h00086;
               12'b010100101111: data1 <=  20'h0e887;
               12'b010100110000: data1 <=  20'h07049;
               12'b010100110001: data1 <=  20'h36466;
               12'b010100110010: data1 <=  20'h33066;
               12'b010100110011: data1 <=  20'h428a5;
               12'b010100110100: data1 <=  20'h3f4a5;
               12'b010100110101: data1 <=  20'h304c3;
               12'b010100110110: data1 <=  20'h4b4c5;
               12'b010100110111: data1 <=  20'h620c4;
               12'b010100111000: data1 <=  20'h0c982;
               12'b010100111001: data1 <=  20'h0a033;
               12'b010100111010: data1 <=  20'h08433;
               12'b010100111011: data1 <=  20'h0bc34;
               12'b010100111100: data1 <=  20'h06834;
               12'b010100111101: data1 <=  20'h49c4c;
               12'b010100111110: data1 <=  20'h4544c;
               12'b010100111111: data1 <=  20'h52247;
               12'b010101000000: data1 <=  20'h590e4;
               12'b010101000001: data1 <=  20'h53184;
               12'b010101000010: data1 <=  20'h73525;
               12'b010101000011: data1 <=  20'h8aa81;
               12'b010101000100: data1 <=  20'h4d466;
               12'b010101000101: data1 <=  20'h2ce41;
               12'b010101000110: data1 <=  20'h2ca41;
               12'b010101000111: data1 <=  20'h304c3;
               12'b010101001000: data1 <=  20'h58122;
               12'b010101001001: data1 <=  20'h5ad22;
               12'b010101001010: data1 <=  20'h2d867;
               12'b010101001011: data1 <=  20'h548c3;
               12'b010101001100: data1 <=  20'h2e489;
               12'b010101001101: data1 <=  20'h4e066;
               12'b010101001110: data1 <=  20'h2bc85;
               12'b010101001111: data1 <=  20'h02c66;
               12'b010101010000: data1 <=  20'h4b983;
               12'b010101010001: data1 <=  20'h548c3;
               12'b010101010010: data1 <=  20'h528c3;
               12'b010101010011: data1 <=  20'h6c922;
               12'b010101010100: data1 <=  20'h78183;
               12'b010101010101: data1 <=  20'h13a81;
               12'b010101010110: data1 <=  20'h20c86;
               12'b010101010111: data1 <=  20'h03038;
               12'b010101011000: data1 <=  20'h660a4;
               12'b010101011001: data1 <=  20'h72cc6;
               12'b010101011010: data1 <=  20'h5e0c4;
               12'b010101011011: data1 <=  20'h43487;
               12'b010101011100: data1 <=  20'h38887;
               12'b010101011101: data1 <=  20'h66525;
               12'b010101011110: data1 <=  20'h39d82;
               12'b010101011111: data1 <=  20'h60c49;
               12'b010101100000: data1 <=  20'h34867;
               12'b010101100001: data1 <=  20'h1c885;
               12'b010101100010: data1 <=  20'h394c3;
               12'b010101100011: data1 <=  20'h2790c;
               12'b010101100100: data1 <=  20'h2d46e;
               12'b010101100101: data1 <=  20'h4fca4;
               12'b010101100110: data1 <=  20'h4b0a4;
               12'b010101100111: data1 <=  20'h29cc3;
               12'b010101101000: data1 <=  20'h25cc3;
               12'b010101101001: data1 <=  20'h23cc3;
               12'b010101101010: data1 <=  20'h1f4c3;
               12'b010101101011: data1 <=  20'h20242;
               12'b010101101100: data1 <=  20'h1fd22;
               12'b010101101101: data1 <=  20'h164a4;
               12'b010101101110: data1 <=  20'h140a4;
               12'b010101101111: data1 <=  20'h4746c;
               12'b010101110000: data1 <=  20'h4786b;
               12'b010101110001: data1 <=  20'h33ca4;
               12'b010101110010: data1 <=  20'h28867;
               12'b010101110011: data1 <=  20'h78241;
               12'b010101110100: data1 <=  20'h1b849;
               12'b010101110101: data1 <=  20'h09067;
               12'b010101110110: data1 <=  20'h47066;
               12'b010101110111: data1 <=  20'h4e84b;
               12'b010101111000: data1 <=  20'h4d04b;
               12'b010101111001: data1 <=  20'h03092;
               12'b010101111010: data1 <=  20'h4cca5;
               12'b010101111011: data1 <=  20'h83ec1;
               12'b010101111100: data1 <=  20'h19434;
               12'b010101111101: data1 <=  20'h0e904;
               12'b010101111110: data1 <=  20'h40542;
               12'b010101111111: data1 <=  20'h2d485;
               12'b010110000000: data1 <=  20'h04467;
               12'b010110000001: data1 <=  20'h5eca4;
               12'b010110000010: data1 <=  20'h13683;
               12'b010110000011: data1 <=  20'h2d4c4;
               12'b010110000100: data1 <=  20'h7f4c3;
               12'b010110000101: data1 <=  20'h4cd42;
               12'b010110000110: data1 <=  20'h21c89;
               12'b010110000111: data1 <=  20'h46c68;
               12'b010110001000: data1 <=  20'h1d851;
               12'b010110001001: data1 <=  20'h00c66;
               12'b010110001010: data1 <=  20'h1d851;
               12'b010110001011: data1 <=  20'h1a051;
               12'b010110001100: data1 <=  20'h78261;
               12'b010110001101: data1 <=  20'h3b049;
               12'b010110001110: data1 <=  20'h55049;
               12'b010110001111: data1 <=  20'h53049;
               12'b010110010000: data1 <=  20'h47ca4;
               12'b010110010001: data1 <=  20'h28849;
               12'b010110010010: data1 <=  20'h03049;
               12'b010110010011: data1 <=  20'h38d04;
               12'b010110010100: data1 <=  20'h740c3;
               12'b010110010101: data1 <=  20'h2e449;
               12'b010110010110: data1 <=  20'h740c3;
               12'b010110010111: data1 <=  20'h58582;
               12'b010110011000: data1 <=  20'h5b122;
               12'b010110011001: data1 <=  20'h57d22;
               12'b010110011010: data1 <=  20'h32e41;
               12'b010110011011: data1 <=  20'h38ac2;
               12'b010110011100: data1 <=  20'h304c3;
               12'b010110011101: data1 <=  20'h2bcc3;
               12'b010110011110: data1 <=  20'h58e03;
               12'b010110011111: data1 <=  20'h72122;
               12'b010110100000: data1 <=  20'h740c3;
               12'b010110100001: data1 <=  20'h718c3;
               12'b010110100010: data1 <=  20'h0a857;
               12'b010110100011: data1 <=  20'h85503;
               12'b010110100100: data1 <=  20'h7f104;
               12'b010110100101: data1 <=  20'h07857;
               12'b010110100110: data1 <=  20'h71641;
               12'b010110100111: data1 <=  20'h6a641;
               12'b010110101000: data1 <=  20'h67162;
               12'b010110101001: data1 <=  20'h70922;
               12'b010110101010: data1 <=  20'h40ce3;
               12'b010110101011: data1 <=  20'h710c3;
               12'b010110101100: data1 <=  20'h2bf02;
               12'b010110101101: data1 <=  20'h2e485;
               12'b010110101110: data1 <=  20'h53cc6;
               12'b010110101111: data1 <=  20'h27849;
               12'b010110110000: data1 <=  20'h03449;
               12'b010110110001: data1 <=  20'h2e849;
               12'b010110110010: data1 <=  20'h0d281;
               12'b010110110011: data1 <=  20'h70cc3;
               12'b010110110100: data1 <=  20'h0fc4d;
               12'b010110110101: data1 <=  20'h2ecc4;
               12'b010110110110: data1 <=  20'h08c4d;
               12'b010110110111: data1 <=  20'h01c32;
               12'b010110111000: data1 <=  20'h164a5;
               12'b010110111001: data1 <=  20'h60488;
               12'b010110111010: data1 <=  20'h41449;
               12'b010110111011: data1 <=  20'h15449;
               12'b010110111100: data1 <=  20'h05067;
               12'b010110111101: data1 <=  20'h00467;
               12'b010110111110: data1 <=  20'h04468;
               12'b010110111111: data1 <=  20'h1b44a;
               12'b010111000000: data1 <=  20'h6d523;
               12'b010111000001: data1 <=  20'h80164;
               12'b010111000010: data1 <=  20'h164a5;
               12'b010111000011: data1 <=  20'h140a5;
               12'b010111000100: data1 <=  20'h29890;
               12'b010111000101: data1 <=  20'h26890;
               12'b010111000110: data1 <=  20'h5a0a5;
               12'b010111000111: data1 <=  20'h772a1;
               12'b010111001000: data1 <=  20'h10522;
               12'b010111001001: data1 <=  20'h094c4;
               12'b010111001010: data1 <=  20'h030c6;
               12'b010111001011: data1 <=  20'h40886;
               12'b010111001100: data1 <=  20'h68ca4;
               12'b010111001101: data1 <=  20'h640a4;
               12'b010111001110: data1 <=  20'h4e885;
               12'b010111001111: data1 <=  20'h658a4;
               12'b010111010000: data1 <=  20'h28cc3;
               12'b010111010001: data1 <=  20'h27c49;
               12'b010111010010: data1 <=  20'h3b867;
               12'b010111010011: data1 <=  20'h3a467;
               12'b010111010100: data1 <=  20'h40566;
               12'b010111010101: data1 <=  20'h33068;
               12'b010111010110: data1 <=  20'h42c87;
               12'b010111010111: data1 <=  20'h3f487;
               12'b010111011000: data1 <=  20'h09c89;
               12'b010111011001: data1 <=  20'h1fd04;
               12'b010111011010: data1 <=  20'h3f644;
               12'b010111011011: data1 <=  20'h58a04;
               12'b010111011100: data1 <=  20'h1dc8a;
               12'b010111011101: data1 <=  20'h0f066;
               12'b010111011110: data1 <=  20'h1dc8a;
               12'b010111011111: data1 <=  20'h1948a;
               12'b010111100000: data1 <=  20'h35c87;
               12'b010111100001: data1 <=  20'h33487;
               12'b010111100010: data1 <=  20'h6cca4;
               12'b010111100011: data1 <=  20'h650e3;
               12'b010111100100: data1 <=  20'h70b05;
               12'b010111100101: data1 <=  20'h0e88b;
               12'b010111100110: data1 <=  20'h10088;
               12'b010111100111: data1 <=  20'h0c983;
               12'b010111101000: data1 <=  20'h14583;
               12'b010111101001: data1 <=  20'h0ccc6;
               12'b010111101010: data1 <=  20'h368c3;
               12'b010111101011: data1 <=  20'h13c85;
               12'b010111101100: data1 <=  20'h8b241;
               12'b010111101101: data1 <=  20'h45241;
               12'b010111101110: data1 <=  20'h452c1;
               12'b010111101111: data1 <=  20'h45583;
               12'b010111110000: data1 <=  20'h368c3;
               12'b010111110001: data1 <=  20'h320c3;
               12'b010111110010: data1 <=  20'h60c49;
               12'b010111110011: data1 <=  20'h5f922;
               12'b010111110100: data1 <=  20'h59ce6;
               12'b010111110101: data1 <=  20'h53066;
               12'b010111110110: data1 <=  20'h60cc4;
               12'b010111110111: data1 <=  20'h1ac50;
               12'b010111111000: data1 <=  20'h60c49;
               12'b010111111001: data1 <=  20'h60449;
               12'b010111111010: data1 <=  20'h488c5;
               12'b010111111011: data1 <=  20'h32dc2;
               12'b010111111100: data1 <=  20'h26a24;
               12'b010111111101: data1 <=  20'h39d87;
               12'b010111111110: data1 <=  20'h1b123;
               12'b010111111111: data1 <=  20'h2ed83;
               12'b011000000000: data1 <=  20'h47925;
               12'b011000000001: data1 <=  20'h4ba41;
               12'b011000000010: data1 <=  20'h72922;
               12'b011000000011: data1 <=  20'h0c922;
               12'b011000000100: data1 <=  20'h51702;
               12'b011000000101: data1 <=  20'h4ba83;
               12'b011000000110: data1 <=  20'h22506;
               12'b011000000111: data1 <=  20'h2e485;
               12'b011000001000: data1 <=  20'h21142;
               12'b011000001001: data1 <=  20'h790c4;
               12'b011000001010: data1 <=  20'h238e5;
               12'b011000001011: data1 <=  20'h1f4e5;
               12'b011000001100: data1 <=  20'h0b066;
               12'b011000001101: data1 <=  20'h19664;
               12'b011000001110: data1 <=  20'h1c122;
               12'b011000001111: data1 <=  20'h19d22;
               12'b011000010000: data1 <=  20'h1c142;
               12'b011000010001: data1 <=  20'h1c122;
               12'b011000010010: data1 <=  20'h09449;
               12'b011000010011: data1 <=  20'h08c49;
               12'b011000010100: data1 <=  20'h22c85;
               12'b011000010101: data1 <=  20'h1b88d;
               12'b011000010110: data1 <=  20'h22866;
               12'b011000010111: data1 <=  20'h210c3;
               12'b011000011000: data1 <=  20'h2d942;
               12'b011000011001: data1 <=  20'h024e5;
               12'b011000011010: data1 <=  20'h44d23;
               12'b011000011011: data1 <=  20'h28449;
               12'b011000011100: data1 <=  20'h13867;
               12'b011000011101: data1 <=  20'h744c3;
               12'b011000011110: data1 <=  20'h32943;
               12'b011000011111: data1 <=  20'h1c542;
               12'b011000100000: data1 <=  20'h45ca6;
               12'b011000100001: data1 <=  20'h1e049;
               12'b011000100010: data1 <=  20'h53507;
               12'b011000100011: data1 <=  20'h09583;
               12'b011000100100: data1 <=  20'h19849;
               12'b011000100101: data1 <=  20'h2ca41;
               12'b011000100110: data1 <=  20'h77a02;
               12'b011000100111: data1 <=  20'h3b8c3;
               12'b011000101000: data1 <=  20'h26ce3;
               12'b011000101001: data1 <=  20'h23885;
               12'b011000101010: data1 <=  20'h13681;
               12'b011000101011: data1 <=  20'h0f866;
               12'b011000101100: data1 <=  20'h28049;
               12'b011000101101: data1 <=  20'h15c4b;
               12'b011000101110: data1 <=  20'h1544b;
               12'b011000101111: data1 <=  20'h15c85;
               12'b011000110000: data1 <=  20'h09432;
               12'b011000110001: data1 <=  20'h0f866;
               12'b011000110010: data1 <=  20'h12e61;
               12'b011000110011: data1 <=  20'h66522;
               12'b011000110100: data1 <=  20'h33cc5;
               12'b011000110101: data1 <=  20'h03849;
               12'b011000110110: data1 <=  20'h02049;
               12'b011000110111: data1 <=  20'h48085;
               12'b011000111000: data1 <=  20'h25e41;
               12'b011000111001: data1 <=  20'h3a9c2;
               12'b011000111010: data1 <=  20'h6ae41;
               12'b011000111011: data1 <=  20'h7a922;
               12'b011000111100: data1 <=  20'h320c3;
               12'b011000111101: data1 <=  20'h6c8e4;
               12'b011000111110: data1 <=  20'h71281;
               12'b011000111111: data1 <=  20'h7a922;
               12'b011001000000: data1 <=  20'h0d9e2;
               12'b011001000001: data1 <=  20'h238c3;
               12'b011001000010: data1 <=  20'h258c3;
               12'b011001000011: data1 <=  20'h7a922;
               12'b011001000100: data1 <=  20'h76d22;
               12'b011001000101: data1 <=  20'h744c3;
               12'b011001000110: data1 <=  20'h714c3;
               12'b011001000111: data1 <=  20'h56485;
               12'b011001001000: data1 <=  20'h59904;
               12'b011001001001: data1 <=  20'h73c66;
               12'b011001001010: data1 <=  20'h51485;
               12'b011001001011: data1 <=  20'h6a703;
               12'b011001001100: data1 <=  20'h0dcc4;
               12'b011001001101: data1 <=  20'h3b066;
               12'b011001001110: data1 <=  20'h20602;
               12'b011001001111: data1 <=  20'h2e485;
               12'b011001010000: data1 <=  20'h340a4;
               12'b011001010001: data1 <=  20'h3b124;
               12'b011001010010: data1 <=  20'h39524;
               12'b011001010011: data1 <=  20'h3bcc3;
               12'b011001010100: data1 <=  20'h32a84;
               12'b011001010101: data1 <=  20'h4c228;
               12'b011001010110: data1 <=  20'h408e3;
               12'b011001010111: data1 <=  20'h3eee1;
               12'b011001011000: data1 <=  20'h02449;
               12'b011001011001: data1 <=  20'h16049;
               12'b011001011010: data1 <=  20'h08c4d;
               12'b011001011011: data1 <=  20'h90e41;
               12'b011001011100: data1 <=  20'h40066;
               12'b011001011101: data1 <=  20'h03838;
               12'b011001011110: data1 <=  20'h02438;
               12'b011001011111: data1 <=  20'h0ecca;
               12'b011001100000: data1 <=  20'h538a6;
               12'b011001100001: data1 <=  20'h858c3;
               12'b011001100010: data1 <=  20'h0904b;
               12'b011001100011: data1 <=  20'h2e0a4;
               12'b011001100100: data1 <=  20'h030b2;
               12'b011001100101: data1 <=  20'h09c50;
               12'b011001100110: data1 <=  20'h08450;
               12'b011001100111: data1 <=  20'h23cc3;
               12'b011001101000: data1 <=  20'h26641;
               12'b011001101001: data1 <=  20'h23cc3;
               12'b011001101010: data1 <=  20'h1f4c3;
               12'b011001101011: data1 <=  20'h54962;
               12'b011001101100: data1 <=  20'h2e4a4;
               12'b011001101101: data1 <=  20'h3b0a7;
               12'b011001101110: data1 <=  20'h3a4a7;
               12'b011001101111: data1 <=  20'h1d066;
               12'b011001110000: data1 <=  20'h26ca4;
               12'b011001110001: data1 <=  20'h85103;
               12'b011001110010: data1 <=  20'h85903;
               12'b011001110011: data1 <=  20'h22967;
               12'b011001110100: data1 <=  20'h3f485;
               12'b011001110101: data1 <=  20'h05066;
               12'b011001110110: data1 <=  20'h0e452;
               12'b011001110111: data1 <=  20'h03c49;
               12'b011001111000: data1 <=  20'h5dce3;
               12'b011001111001: data1 <=  20'h56085;
               12'b011001111010: data1 <=  20'h00466;
               12'b011001111011: data1 <=  20'h2ec66;
               12'b011001111100: data1 <=  20'h51885;
               12'b011001111101: data1 <=  20'h8a661;
               12'b011001111110: data1 <=  20'h14c4d;
               12'b011001111111: data1 <=  20'h46241;
               12'b011010000000: data1 <=  20'h2e0a4;
               12'b011010000001: data1 <=  20'h2e885;
               12'b011010000010: data1 <=  20'h13e02;
               12'b011010000011: data1 <=  20'h07e41;
               12'b011010000100: data1 <=  20'h078a4;
               12'b011010000101: data1 <=  20'h74cc3;
               12'b011010000110: data1 <=  20'h608c3;
               12'b011010000111: data1 <=  20'h3ed64;
               12'b011010001000: data1 <=  20'h3ac66;
               12'b011010001001: data1 <=  20'h47485;
               12'b011010001010: data1 <=  20'h2e8a7;
               12'b011010001011: data1 <=  20'h0f48a;
               12'b011010001100: data1 <=  20'h0ec8a;
               12'b011010001101: data1 <=  20'h1cd23;
               12'b011010001110: data1 <=  20'h32143;
               12'b011010001111: data1 <=  20'h38ea2;
               12'b011010010000: data1 <=  20'h19168;
               12'b011010010001: data1 <=  20'h470cb;
               12'b011010010010: data1 <=  20'h2e066;
               12'b011010010011: data1 <=  20'h048c9;
               12'b011010010100: data1 <=  20'h000c9;
               12'b011010010101: data1 <=  20'h09562;
               12'b011010010110: data1 <=  20'h0d642;
               12'b011010010111: data1 <=  20'h2c6c2;
               12'b011010011000: data1 <=  20'h140c3;
               12'b011010011001: data1 <=  20'h5a849;
               12'b011010011010: data1 <=  20'h5a049;
               12'b011010011011: data1 <=  20'h78241;
               12'b011010011100: data1 <=  20'h0246d;
               12'b011010011101: data1 <=  20'h1acc4;
               12'b011010011110: data1 <=  20'h0ec86;
               12'b011010011111: data1 <=  20'h0da41;
               12'b011010100000: data1 <=  20'h4b0c4;
               12'b011010100001: data1 <=  20'h60849;
               12'b011010100010: data1 <=  20'h4144d;
               12'b011010100011: data1 <=  20'h72241;
               12'b011010100100: data1 <=  20'h1bc49;
               12'b011010100101: data1 <=  20'h03049;
               12'b011010100110: data1 <=  20'h26ca4;
               12'b011010100111: data1 <=  20'h54ca4;
               12'b011010101000: data1 <=  20'h528a4;
               12'b011010101001: data1 <=  20'h54d22;
               12'b011010101010: data1 <=  20'h2bee5;
               12'b011010101011: data1 <=  20'h29906;
               12'b011010101100: data1 <=  20'h718c3;
               12'b011010101101: data1 <=  20'h7f122;
               12'b011010101110: data1 <=  20'h70a41;
               12'b011010101111: data1 <=  20'h54962;
               12'b011010110000: data1 <=  20'h51562;
               12'b011010110001: data1 <=  20'h3b583;
               12'b011010110010: data1 <=  20'h7e904;
               12'b011010110011: data1 <=  20'h731c2;
               12'b011010110100: data1 <=  20'h0cea1;
               12'b011010110101: data1 <=  20'h0c983;
               12'b011010110110: data1 <=  20'h5f485;
               12'b011010110111: data1 <=  20'h470e3;
               12'b011010111000: data1 <=  20'h70cc3;
               12'b011010111001: data1 <=  20'h79485;
               12'b011010111010: data1 <=  20'h4cc85;
               12'b011010111011: data1 <=  20'h4d4c4;
               12'b011010111100: data1 <=  20'h08c66;
               12'b011010111101: data1 <=  20'h5ea61;
               12'b011010111110: data1 <=  20'h2d8a5;
               12'b011010111111: data1 <=  20'h4bd2c;
               12'b011011000000: data1 <=  20'h0284c;
               12'b011011000001: data1 <=  20'h13a23;
               12'b011011000010: data1 <=  20'h0288b;
               12'b011011000011: data1 <=  20'h0106d;
               12'b011011000100: data1 <=  20'h46203;
               12'b011011000101: data1 <=  20'h598a6;
               12'b011011000110: data1 <=  20'h858c3;
               12'b011011000111: data1 <=  20'h00c66;
               12'b011011001000: data1 <=  20'h06e81;
               12'b011011001001: data1 <=  20'h27caa;
               12'b011011001010: data1 <=  20'h28449;
               12'b011011001011: data1 <=  20'h02c49;
               12'b011011001100: data1 <=  20'h04049;
               12'b011011001101: data1 <=  20'h72522;
               12'b011011001110: data1 <=  20'h04049;
               12'b011011001111: data1 <=  20'h01849;
               12'b011011010000: data1 <=  20'h0b050;
               12'b011011010001: data1 <=  20'h07050;
               12'b011011010010: data1 <=  20'h678c3;
               12'b011011010011: data1 <=  20'h12cc3;
               12'b011011010100: data1 <=  20'h21866;
               12'b011011010101: data1 <=  20'h40066;
               12'b011011010110: data1 <=  20'h61468;
               12'b011011010111: data1 <=  20'h3f8e6;
               12'b011011011000: data1 <=  20'h33d82;
               12'b011011011001: data1 <=  20'h0ec54;
               12'b011011011010: data1 <=  20'h678c3;
               12'b011011011011: data1 <=  20'h28849;
               12'b011011011100: data1 <=  20'h678c3;
               12'b011011011101: data1 <=  20'h8adc2;
               12'b011011011110: data1 <=  20'h3fa06;
               12'b011011011111: data1 <=  20'h28449;
               12'b011011100000: data1 <=  20'h0d6a2;
               12'b011011100001: data1 <=  20'h650c3;
               12'b011011100010: data1 <=  20'h810a4;
               12'b011011100011: data1 <=  20'h01108;
               12'b011011100100: data1 <=  20'h28ce3;
               12'b011011100101: data1 <=  20'h41085;
               12'b011011100110: data1 <=  20'h618c4;
               12'b011011100111: data1 <=  20'h2ecc4;
               12'b011011101000: data1 <=  20'h288e3;
               12'b011011101001: data1 <=  20'h26525;
               12'b011011101010: data1 <=  20'h030d5;
               12'b011011101011: data1 <=  20'h02115;
               12'b011011101100: data1 <=  20'h78641;
               12'b011011101101: data1 <=  20'h6a522;
               12'b011011101110: data1 <=  20'h1a261;
               12'b011011101111: data1 <=  20'h19301;
               12'b011011110000: data1 <=  20'h67d22;
               12'b011011110001: data1 <=  20'h64122;
               12'b011011110010: data1 <=  20'h65a41;
               12'b011011110011: data1 <=  20'h71641;
               12'b011011110100: data1 <=  20'h03437;
               12'b011011110101: data1 <=  20'h14503;
               12'b011011110110: data1 <=  20'h6be41;
               12'b011011110111: data1 <=  20'h02837;
               12'b011011111000: data1 <=  20'h4d885;
               12'b011011111001: data1 <=  20'h4cd44;
               12'b011011111010: data1 <=  20'h3c867;
               12'b011011111011: data1 <=  20'h13543;
               12'b011011111100: data1 <=  20'h2e8a6;
               12'b011011111101: data1 <=  20'h194c5;
               12'b011011111110: data1 <=  20'h16922;
               12'b011011111111: data1 <=  20'h0cc85;
               12'b011100000000: data1 <=  20'h21ca4;
               12'b011100000001: data1 <=  20'h02cf8;
               12'b011100000010: data1 <=  20'h78942;
               12'b011100000011: data1 <=  20'h79485;
               12'b011100000100: data1 <=  20'h61849;
               12'b011100000101: data1 <=  20'h8a641;
               12'b011100000110: data1 <=  20'h61849;
               12'b011100000111: data1 <=  20'h5f849;
               12'b011100001000: data1 <=  20'h28849;
               12'b011100001001: data1 <=  20'h1504b;
               12'b011100001010: data1 <=  20'h16922;
               12'b011100001011: data1 <=  20'h335c4;
               12'b011100001100: data1 <=  20'h1b1e3;
               12'b011100001101: data1 <=  20'h0e485;
               12'b011100001110: data1 <=  20'h0f86c;
               12'b011100001111: data1 <=  20'h0ec6c;
               12'b011100010000: data1 <=  20'h2d8c4;
               12'b011100010001: data1 <=  20'h1548a;
               12'b011100010010: data1 <=  20'h28d03;
               12'b011100010011: data1 <=  20'h088c9;
               12'b011100010100: data1 <=  20'h344c5;
               12'b011100010101: data1 <=  20'h0018b;
               12'b011100010110: data1 <=  20'h74122;
               12'b011100010111: data1 <=  20'h7d304;
               12'b011100011000: data1 <=  20'h79d62;
               12'b011100011001: data1 <=  20'h70d22;
               12'b011100011010: data1 <=  20'h33ca4;
               12'b011100011011: data1 <=  20'h60849;
               12'b011100011100: data1 <=  20'h748c3;
               12'b011100011101: data1 <=  20'h710c3;
               12'b011100011110: data1 <=  20'h27a03;
               12'b011100011111: data1 <=  20'h2bd42;
               12'b011100100000: data1 <=  20'h26e41;
               12'b011100100001: data1 <=  20'h38d23;
               12'b011100100010: data1 <=  20'h22d43;
               12'b011100100011: data1 <=  20'h2ca41;
               12'b011100100100: data1 <=  20'h1b5e2;
               12'b011100100101: data1 <=  20'h3f9e2;
               12'b011100100110: data1 <=  20'h22582;
               12'b011100100111: data1 <=  20'h3444c;
               12'b011100101000: data1 <=  20'h03449;
               12'b011100101001: data1 <=  20'h4b066;
               12'b011100101010: data1 <=  20'h5b142;
               12'b011100101011: data1 <=  20'h3f243;
               12'b011100101100: data1 <=  20'h6d143;
               12'b011100101101: data1 <=  20'h274a4;
               12'b011100101110: data1 <=  20'h28ce3;
               12'b011100101111: data1 <=  20'h53067;
               12'b011100110000: data1 <=  20'h42c66;
               12'b011100110001: data1 <=  20'h3f866;
               12'b011100110010: data1 <=  20'h3b886;
               12'b011100110011: data1 <=  20'h1544e;
               12'b011100110100: data1 <=  20'h04832;
               12'b011100110101: data1 <=  20'h4e10c;
               12'b011100110110: data1 <=  20'h0444e;
               12'b011100110111: data1 <=  20'h0144e;
               12'b011100111000: data1 <=  20'h10894;
               12'b011100111001: data1 <=  20'h0d894;
               12'b011100111010: data1 <=  20'h04851;
               12'b011100111011: data1 <=  20'h01051;
               12'b011100111100: data1 <=  20'h35d22;
               12'b011100111101: data1 <=  20'h32122;
               12'b011100111110: data1 <=  20'h0b44d;
               12'b011100111111: data1 <=  20'h06c4d;
               12'b011101000000: data1 <=  20'h04049;
               12'b011101000001: data1 <=  20'h40c87;
               12'b011101000010: data1 <=  20'h47d82;
               12'b011101000011: data1 <=  20'h44d82;
               12'b011101000100: data1 <=  20'h3fdc3;
               12'b011101000101: data1 <=  20'h64281;
               12'b011101000110: data1 <=  20'h41885;
               12'b011101000111: data1 <=  20'h2d1a3;
               12'b011101001000: data1 <=  20'h348c6;
               12'b011101001001: data1 <=  20'h02049;
               12'b011101001010: data1 <=  20'h46582;
               12'b011101001011: data1 <=  20'h265e4;
               12'b011101001100: data1 <=  20'h04085;
               12'b011101001101: data1 <=  20'h5f4c3;
               12'b011101001110: data1 <=  20'h59905;
               12'b011101001111: data1 <=  20'h07c32;
               12'b011101010000: data1 <=  20'h0284e;
               12'b011101010001: data1 <=  20'h15849;
               12'b011101010010: data1 <=  20'h100c3;
               12'b011101010011: data1 <=  20'h25a22;
               12'b011101010100: data1 <=  20'h810a4;
               12'b011101010101: data1 <=  20'h7dca4;
               12'b011101010110: data1 <=  20'h78641;
               12'b011101010111: data1 <=  20'h01085;
               12'b011101011000: data1 <=  20'h17066;
               12'b011101011001: data1 <=  20'h4b84c;
               12'b011101011010: data1 <=  20'h19aa1;
               12'b011101011011: data1 <=  20'h13c66;
               12'b011101011100: data1 <=  20'h368c3;
               12'b011101011101: data1 <=  20'h5fd09;
               12'b011101011110: data1 <=  20'h52d25;
               12'b011101011111: data1 <=  20'h270a6;
               12'b011101100000: data1 <=  20'h3bc66;
               12'b011101100001: data1 <=  20'h020ab;
               12'b011101100010: data1 <=  20'h3c066;
               12'b011101100011: data1 <=  20'h39c66;
               12'b011101100100: data1 <=  20'h22ca4;
               12'b011101100101: data1 <=  20'h1a104;
               12'b011101100110: data1 <=  20'h2d8c3;
               12'b011101100111: data1 <=  20'h0206d;
               12'b011101101000: data1 <=  20'h03449;
               12'b011101101001: data1 <=  20'h02449;
               12'b011101101010: data1 <=  20'h1b143;
               12'b011101101011: data1 <=  20'h12e41;
               12'b011101101100: data1 <=  20'h558e3;
               12'b011101101101: data1 <=  20'h514e3;
               12'b011101101110: data1 <=  20'h11c35;
               12'b011101101111: data1 <=  20'h514a4;
               12'b011101110000: data1 <=  20'h35182;
               12'b011101110001: data1 <=  20'h38a81;
               12'b011101110010: data1 <=  20'h33661;
               12'b011101110011: data1 <=  20'h57d22;
               12'b011101110100: data1 <=  20'h591c4;
               12'b011101110101: data1 <=  20'h4c5c6;
               12'b011101110110: data1 <=  20'h4e867;
               12'b011101110111: data1 <=  20'h6aa42;
               12'b011101111000: data1 <=  20'h6d0c3;
               12'b011101111001: data1 <=  20'h32122;
               12'b011101111010: data1 <=  20'h41d43;
               12'b011101111011: data1 <=  20'h3ed43;
               12'b011101111100: data1 <=  20'h38582;
               12'b011101111101: data1 <=  20'h4b544;
               12'b011101111110: data1 <=  20'h4e867;
               12'b011101111111: data1 <=  20'h4cc67;
               12'b011110000000: data1 <=  20'h4e085;
               12'b011110000001: data1 <=  20'h4d085;
               12'b011110000010: data1 <=  20'h41c4a;
               12'b011110000011: data1 <=  20'h60942;
               12'b011110000100: data1 <=  20'h40c66;
               12'b011110000101: data1 <=  20'h080e3;
               12'b011110000110: data1 <=  20'h2d5a3;
               12'b011110000111: data1 <=  20'h21c85;
               12'b011110001000: data1 <=  20'h4d942;
               12'b011110001001: data1 <=  20'h658a4;
               12'b011110001010: data1 <=  20'h03c49;
               12'b011110001011: data1 <=  20'h408c6;
               12'b011110001100: data1 <=  20'h1bd22;
               12'b011110001101: data1 <=  20'h7f0e3;
               12'b011110001110: data1 <=  20'h452c1;
               12'b011110001111: data1 <=  20'h70a41;
               12'b011110010000: data1 <=  20'h03c49;
               12'b011110010001: data1 <=  20'h01c49;
               12'b011110010010: data1 <=  20'h11854;
               12'b011110010011: data1 <=  20'h0d054;
               12'b011110010100: data1 <=  20'h2f467;
               12'b011110010101: data1 <=  20'h06c49;
               12'b011110010110: data1 <=  20'h67122;
               12'b011110010111: data1 <=  20'h5e122;
               12'b011110011000: data1 <=  20'h33de2;
               12'b011110011001: data1 <=  20'h34066;
               12'b011110011010: data1 <=  20'h288c3;
               12'b011110011011: data1 <=  20'h77542;
               12'b011110011100: data1 <=  20'h740c3;
               12'b011110011101: data1 <=  20'h20127;
               12'b011110011110: data1 <=  20'h29c49;
               12'b011110011111: data1 <=  20'h26c49;
               12'b011110100000: data1 <=  20'h03449;
               12'b011110100001: data1 <=  20'h02449;
               12'b011110100010: data1 <=  20'h22849;
               12'b011110100011: data1 <=  20'h22466;
               12'b011110100100: data1 <=  20'h09503;
               12'b011110100101: data1 <=  20'h5404b;
               12'b011110100110: data1 <=  20'h0b466;
               12'b011110100111: data1 <=  20'h70e41;
               12'b011110101000: data1 <=  20'h6c144;
               12'b011110101001: data1 <=  20'h7e942;
               12'b011110101010: data1 <=  20'h66522;
               12'b011110101011: data1 <=  20'h06866;
               12'b011110101100: data1 <=  20'h36ca4;
               12'b011110101101: data1 <=  20'h01088;
               12'b011110101110: data1 <=  20'h26661;
               12'b011110101111: data1 <=  20'h1f8c3;
               12'b011110110000: data1 <=  20'h088e8;
               12'b011110110001: data1 <=  20'h20604;
               12'b011110110010: data1 <=  20'h07e41;
               12'b011110110011: data1 <=  20'h45d47;
               12'b011110110100: data1 <=  20'h48885;
               12'b011110110101: data1 <=  20'h72cc3;
               12'b011110110110: data1 <=  20'h73886;
               12'b011110110111: data1 <=  20'h5f469;
               12'b011110111000: data1 <=  20'h488c4;
               12'b011110111001: data1 <=  20'h458c4;
               12'b011110111010: data1 <=  20'h3bd23;
               12'b011110111011: data1 <=  20'h5e182;
               12'b011110111100: data1 <=  20'h6dd42;
               12'b011110111101: data1 <=  20'h6a542;
               12'b011110111110: data1 <=  20'h67cc3;
               12'b011110111111: data1 <=  20'h64cc3;
               12'b011111000000: data1 <=  20'h21888;
               12'b011111000001: data1 <=  20'h70cc3;
               12'b011111000010: data1 <=  20'h86942;
               12'b011111000011: data1 <=  20'h83942;
               12'b011111000100: data1 <=  20'h7ea41;
               12'b011111000101: data1 <=  20'h78c85;
               12'b011111000110: data1 <=  20'h0cb02;
               12'b011111000111: data1 <=  20'h190c3;
               12'b011111001000: data1 <=  20'h3bd43;
               12'b011111001001: data1 <=  20'h77264;
               12'b011111001010: data1 <=  20'h10142;
               12'b011111001011: data1 <=  20'h408ee;
               12'b011111001100: data1 <=  20'h41088;
               12'b011111001101: data1 <=  20'h34ca4;
               12'b011111001110: data1 <=  20'h21c49;
               12'b011111001111: data1 <=  20'h2184a;
               12'b011111010000: data1 <=  20'h1c84d;
               12'b011111010001: data1 <=  20'h1b04d;
               12'b011111010010: data1 <=  20'h2e866;
               12'b011111010011: data1 <=  20'h26503;
               12'b011111010100: data1 <=  20'h1c507;
               12'b011111010101: data1 <=  20'h00182;
               12'b011111010110: data1 <=  20'h09466;
               12'b011111010111: data1 <=  20'h090e4;
               12'b011111011000: data1 <=  20'h6cce3;
               12'b011111011001: data1 <=  20'h14c85;
               12'b011111011010: data1 <=  20'h15885;
               12'b011111011011: data1 <=  20'h0f04d;
               12'b011111011100: data1 <=  20'h0f833;
               12'b011111011101: data1 <=  20'h2e466;
               12'b011111011110: data1 <=  20'h8a942;
               12'b011111011111: data1 <=  20'h64182;
               12'b011111100000: data1 <=  20'h15885;
               12'b011111100001: data1 <=  20'h3ec87;
               12'b011111100010: data1 <=  20'h798c3;
               12'b011111100011: data1 <=  20'h018ac;
               12'b011111100100: data1 <=  20'h22ce7;
               12'b011111100101: data1 <=  20'h33ca4;
               12'b011111100110: data1 <=  20'h09466;
               12'b011111100111: data1 <=  20'h28983;
               12'b011111101000: data1 <=  20'h15885;
               12'b011111101001: data1 <=  20'h51962;
               12'b011111101010: data1 <=  20'h59d82;
               12'b011111101011: data1 <=  20'h2bd22;
               12'b011111101100: data1 <=  20'h2c2e2;
               12'b011111101101: data1 <=  20'h3ee64;
               12'b011111101110: data1 <=  20'h344c7;
               12'b011111101111: data1 <=  20'h790c3;
               12'b011111110000: data1 <=  20'h5a449;
               12'b011111110001: data1 <=  20'h2844c;
               12'b011111110010: data1 <=  20'h04849;
               12'b011111110011: data1 <=  20'h01049;
               12'b011111110100: data1 <=  20'h0a04b;
               12'b011111110101: data1 <=  20'h57d06;
               12'b011111110110: data1 <=  20'h420e3;
               12'b011111110111: data1 <=  20'h4bd22;
               12'b011111111000: data1 <=  20'h0a04b;
               12'b011111111001: data1 <=  20'h0804b;
               12'b011111111010: data1 <=  20'h2f542;
               12'b011111111011: data1 <=  20'h41867;
               12'b011111111100: data1 <=  20'h2d8a4;
               12'b011111111101: data1 <=  20'h32085;
               12'b011111111110: data1 <=  20'h04c86;
               12'b011111111111: data1 <=  20'h00486;
               12'b100000000000: data1 <=  20'h23450;
               12'b100000000001: data1 <=  20'h20c50;
               12'b100000000010: data1 <=  20'h04450;
               12'b100000000011: data1 <=  20'h01450;
               12'b100000000100: data1 <=  20'h12f01;
               12'b100000000101: data1 <=  20'h14942;
               12'b100000000110: data1 <=  20'h196e4;
               12'b100000000111: data1 <=  20'h70e61;
               12'b100000001000: data1 <=  20'h78641;
               12'b100000001001: data1 <=  20'h77122;
               12'b100000001010: data1 <=  20'h744c3;
               12'b100000001011: data1 <=  20'h714c3;
               12'b100000001100: data1 <=  20'h6b683;
               12'b100000001101: data1 <=  20'h3e867;
               12'b100000001110: data1 <=  20'h78641;
               12'b100000001111: data1 <=  20'h4cc67;
               12'b100000010000: data1 <=  20'h418c5;
               12'b100000010001: data1 <=  20'h400c5;
               12'b100000010010: data1 <=  20'h0ecc9;
               12'b100000010011: data1 <=  20'h268a5;
               12'b100000010100: data1 <=  20'h5c849;
               12'b100000010101: data1 <=  20'h58049;
               12'b100000010110: data1 <=  20'h0984a;
               12'b100000010111: data1 <=  20'h864c3;
               12'b100000011000: data1 <=  20'h0984a;
               12'b100000011001: data1 <=  20'h644a4;
               12'b100000011010: data1 <=  20'h0984a;
               12'b100000011011: data1 <=  20'h00833;
               12'b100000011100: data1 <=  20'h0984a;
               12'b100000011101: data1 <=  20'h06c49;
               12'b100000011110: data1 <=  20'h39262;
               12'b100000011111: data1 <=  20'h65d22;
               12'b100000100000: data1 <=  20'h1d4e3;
               12'b100000100001: data1 <=  20'h1a5c4;
               12'b100000100010: data1 <=  20'h1d103;
               12'b100000100011: data1 <=  20'h19103;
               12'b100000100100: data1 <=  20'h03d22;
               12'b100000100101: data1 <=  20'h64122;
               12'b100000100110: data1 <=  20'h2e0c8;
               12'b100000100111: data1 <=  20'h45c49;
               12'b100000101000: data1 <=  20'h22449;
               12'b100000101001: data1 <=  20'h28049;
               12'b100000101010: data1 <=  20'h0984a;
               12'b100000101011: data1 <=  20'h0884a;
               12'b100000101100: data1 <=  20'h3bd23;
               12'b100000101101: data1 <=  20'h1b049;
               12'b100000101110: data1 <=  20'h66886;
               12'b100000101111: data1 <=  20'h00124;
               12'b100000110000: data1 <=  20'h228e6;
               12'b100000110001: data1 <=  20'h150a7;
               12'b100000110010: data1 <=  20'h5b142;
               12'b100000110011: data1 <=  20'h64085;
               12'b100000110100: data1 <=  20'h452c1;
               12'b100000110101: data1 <=  20'h3ac4a;
               12'b100000110110: data1 <=  20'h10866;
               12'b100000110111: data1 <=  20'h28049;
               12'b100000111000: data1 <=  20'h350a8;
               12'b100000111001: data1 <=  20'h08486;
               12'b100000111010: data1 <=  20'h098c7;
               12'b100000111011: data1 <=  20'h64982;
               12'b100000111100: data1 <=  20'h798c3;
               12'b100000111101: data1 <=  20'h788c3;
               12'b100000111110: data1 <=  20'h1c44a;
               12'b100000111111: data1 <=  20'h7d261;
               12'b100001000000: data1 <=  20'h4e0c4;
               12'b100001000001: data1 <=  20'h4d10b;
               12'b100001000010: data1 <=  20'h4e0c4;
               12'b100001000011: data1 <=  20'h4c8c4;
               12'b100001000100: data1 <=  20'h358c3;
               12'b100001000101: data1 <=  20'h32302;
               12'b100001000110: data1 <=  20'h5b142;
               12'b100001000111: data1 <=  20'h57942;
               12'b100001001000: data1 <=  20'h2ce61;
               12'b100001001001: data1 <=  20'h2c261;
               12'b100001001010: data1 <=  20'h13e03;
               12'b100001001011: data1 <=  20'h08505;
               12'b100001001100: data1 <=  20'h458c5;
               12'b100001001101: data1 <=  20'h28449;
               12'b100001001110: data1 <=  20'h70a41;
               12'b100001001111: data1 <=  20'h91641;
               12'b100001010000: data1 <=  20'h5e4c3;
               12'b100001010001: data1 <=  20'h624c3;
               12'b100001010010: data1 <=  20'h5dcc3;
               12'b100001010011: data1 <=  20'h79885;
               12'b100001010100: data1 <=  20'h59cc8;
               12'b100001010101: data1 <=  20'h4cd45;
               12'b100001010110: data1 <=  20'h1384d;
               12'b100001010111: data1 <=  20'h0ac6d;
               12'b100001011000: data1 <=  20'h08049;
               12'b100001011001: data1 <=  20'h1106b;
               12'b100001011010: data1 <=  20'h0d46b;
               12'b100001011011: data1 <=  20'h59de2;
               12'b100001011100: data1 <=  20'h13681;
               12'b100001011101: data1 <=  20'h28049;
               12'b100001011110: data1 <=  20'h26cc7;
               12'b100001011111: data1 <=  20'h02c49;
               12'b100001100000: data1 <=  20'h02866;
               12'b100001100001: data1 <=  20'h28849;
               12'b100001100010: data1 <=  20'h074ca;
               12'b100001100011: data1 <=  20'h2d523;
               12'b100001100100: data1 <=  20'h2e123;
               12'b100001100101: data1 <=  20'h7f4c3;
               12'b100001100110: data1 <=  20'h28449;
               12'b100001100111: data1 <=  20'h0f08f;
               12'b100001101000: data1 <=  20'h19a41;
               12'b100001101001: data1 <=  20'h1e449;
               12'b100001101010: data1 <=  20'h0ca61;
               12'b100001101011: data1 <=  20'h0dde2;
               12'b100001101100: data1 <=  20'h0f8e5;
               12'b100001101101: data1 <=  20'h0cd6e;
               12'b100001101110: data1 <=  20'h60449;
               12'b100001101111: data1 <=  20'h72241;
               12'b100001110000: data1 <=  20'h4d466;
               12'b100001110001: data1 <=  20'h06e81;
               12'b100001110010: data1 <=  20'h334a4;
               12'b100001110011: data1 <=  20'h28885;
               12'b100001110100: data1 <=  20'h4d466;
               12'b100001110101: data1 <=  20'h5c085;
               12'b100001110110: data1 <=  20'h58085;
               12'b100001110111: data1 <=  20'h748c3;
               12'b100001111000: data1 <=  20'h25cc3;
               12'b100001111001: data1 <=  20'h15c34;
               12'b100001111010: data1 <=  20'h268e3;
               12'b100001111011: data1 <=  20'h21c8d;
               12'b100001111100: data1 <=  20'h39885;
               12'b100001111101: data1 <=  20'h678a4;
               12'b100001111110: data1 <=  20'h33c67;
               12'b100001111111: data1 <=  20'h33d42;
               12'b100010000000: data1 <=  20'h26241;
               12'b100010000001: data1 <=  20'h209e4;
               12'b100010000010: data1 <=  20'h40509;
               12'b100010000011: data1 <=  20'h44f01;
               12'b100010000100: data1 <=  20'h0d04d;
               12'b100010000101: data1 <=  20'h05085;
               12'b100010000110: data1 <=  20'h1a543;
               12'b100010000111: data1 <=  20'h2d241;
               12'b100010001000: data1 <=  20'h0cb01;
               12'b100010001001: data1 <=  20'h1c44b;
               12'b100010001010: data1 <=  20'h00085;
               12'b100010001011: data1 <=  20'h6b641;
               12'b100010001100: data1 <=  20'h6ae41;
               12'b100010001101: data1 <=  20'h03125;
               12'b100010001110: data1 <=  20'h15d55;
               12'b100010001111: data1 <=  20'h2d4e3;
               12'b100010010000: data1 <=  20'h384c3;
               12'b100010010001: data1 <=  20'h5a0e4;
               12'b100010010010: data1 <=  20'h594e4;
               12'b100010010011: data1 <=  20'h860c3;
               12'b100010010100: data1 <=  20'h850c3;
               12'b100010010101: data1 <=  20'h1e449;
               12'b100010010110: data1 <=  20'h32e41;
               12'b100010010111: data1 <=  20'h1e449;
               12'b100010011000: data1 <=  20'h6c142;
               12'b100010011001: data1 <=  20'h66563;
               12'b100010011010: data1 <=  20'h44c85;
               12'b100010011011: data1 <=  20'h74522;
               12'b100010011100: data1 <=  20'h1f849;
               12'b100010011101: data1 <=  20'h35485;
               12'b100010011110: data1 <=  20'h33c85;
               12'b100010011111: data1 <=  20'h35485;
               12'b100010100000: data1 <=  20'h34867;
               12'b100010100001: data1 <=  20'h35485;
               12'b100010100010: data1 <=  20'h28067;
               12'b100010100011: data1 <=  20'h35485;
               12'b100010100100: data1 <=  20'h47486;
               12'b100010100101: data1 <=  20'h461c6;
               12'b100010100110: data1 <=  20'h12d62;
               12'b100010100111: data1 <=  20'h4144a;
               12'b100010101000: data1 <=  20'h77562;
               12'b100010101001: data1 <=  20'h74522;
               12'b100010101010: data1 <=  20'h45241;
               12'b100010101011: data1 <=  20'h1b88d;
               12'b100010101100: data1 <=  20'h76e41;
               12'b100010101101: data1 <=  20'h78641;
               12'b100010101110: data1 <=  20'h70922;
               12'b100010101111: data1 <=  20'h6d922;
               12'b100010110000: data1 <=  20'h6ad22;
               12'b100010110001: data1 <=  20'h09870;
               12'b100010110010: data1 <=  20'h08470;
               12'b100010110011: data1 <=  20'h2284a;
               12'b100010110100: data1 <=  20'h2184a;
               12'b100010110101: data1 <=  20'h03058;
               12'b100010110110: data1 <=  20'h19c4a;
               12'b100010110111: data1 <=  20'h04049;
               12'b100010111000: data1 <=  20'h01849;
               12'b100010111001: data1 <=  20'h21cc5;
               12'b100010111010: data1 <=  20'h27449;
               12'b100010111011: data1 <=  20'h0f8a8;
               12'b100010111100: data1 <=  20'h0e4a8;
               12'b100010111101: data1 <=  20'h02849;
               12'b100010111110: data1 <=  20'h19c66;
               12'b100010111111: data1 <=  20'h04092;
               12'b100011000000: data1 <=  20'h01092;
               12'b100011000001: data1 <=  20'h38702;
               12'b100011000010: data1 <=  20'h2e8e3;
               12'b100011000011: data1 <=  20'h3488f;
               12'b100011000100: data1 <=  20'h030ae;
               12'b100011000101: data1 <=  20'h42c85;
               12'b100011000110: data1 <=  20'h01449;
               12'b100011000111: data1 <=  20'h0a468;
               12'b100011001000: data1 <=  20'h07868;
               12'b100011001001: data1 <=  20'h3f644;
               12'b100011001010: data1 <=  20'h58a02;
               12'b100011001011: data1 <=  20'h58a05;
               12'b100011001100: data1 <=  20'h3f485;
               12'b100011001101: data1 <=  20'h74903;
               12'b100011001110: data1 <=  20'h65885;
               12'b100011001111: data1 <=  20'h67922;
               12'b100011010000: data1 <=  20'h65d22;
               12'b100011010001: data1 <=  20'h58a04;
               12'b100011010010: data1 <=  20'h5de62;
               12'b100011010011: data1 <=  20'h60522;
               12'b100011010100: data1 <=  20'h01837;
               12'b100011010101: data1 <=  20'h3eb02;
               12'b100011010110: data1 <=  20'h384a4;
               12'b100011010111: data1 <=  20'h39269;
               12'b100011011000: data1 <=  20'h47066;
               12'b100011011001: data1 <=  20'h22584;
               12'b100011011010: data1 <=  20'h7e922;
               12'b100011011011: data1 <=  20'h40942;
               12'b100011011100: data1 <=  20'h32a81;
               12'b100011011101: data1 <=  20'h418ea;
               12'b100011011110: data1 <=  20'h3fcea;
               12'b100011011111: data1 <=  20'h48449;
               12'b100011100000: data1 <=  20'h348ac;
               12'b100011100001: data1 <=  20'h3b4c4;
               12'b100011100010: data1 <=  20'h59467;
               12'b100011100011: data1 <=  20'h10cc8;
               12'b100011100100: data1 <=  20'h02449;
               12'b100011100101: data1 <=  20'h67522;
               12'b100011100110: data1 <=  20'h4b162;
               12'b100011100111: data1 <=  20'h4e163;
               12'b100011101000: data1 <=  20'h27c66;
               12'b100011101001: data1 <=  20'h02849;
               12'b100011101010: data1 <=  20'h344c7;
               12'b100011101011: data1 <=  20'h32302;
               12'b100011101100: data1 <=  20'h46d0a;
               12'b100011101101: data1 <=  20'h150d5;
               12'b100011101110: data1 <=  20'h4d44a;
               12'b100011101111: data1 <=  20'h67ca4;
               12'b100011110000: data1 <=  20'h28049;
               12'b100011110001: data1 <=  20'h42466;
               12'b100011110010: data1 <=  20'h40066;
               12'b100011110011: data1 <=  20'h4fc66;
               12'b100011110100: data1 <=  20'h4b866;
               12'b100011110101: data1 <=  20'h60c49;
               12'b100011110110: data1 <=  20'h60449;
               12'b100011110111: data1 <=  20'h808a4;
               12'b100011111000: data1 <=  20'h7e4a4;
               12'b100011111001: data1 <=  20'h79922;
               12'b100011111010: data1 <=  20'h19dc2;
               12'b100011111011: data1 <=  20'h15542;
               12'b100011111100: data1 <=  20'h5f0a4;
               12'b100011111101: data1 <=  20'h11833;
               12'b100011111110: data1 <=  20'h4cc68;
               12'b100011111111: data1 <=  20'h45ca4;
               12'b100100000000: data1 <=  20'h08503;
               12'b100100000001: data1 <=  20'h40182;
               12'b100100000010: data1 <=  20'h1784a;
               12'b100100000011: data1 <=  20'h26466;
               12'b100100000100: data1 <=  20'h05056;
               12'b100100000101: data1 <=  20'h00856;
               12'b100100000110: data1 <=  20'h65661;
               12'b100100000111: data1 <=  20'h4d885;
               12'b100100001000: data1 <=  20'h28449;
               12'b100100001001: data1 <=  20'h89a41;
               12'b100100001010: data1 <=  20'h33d45;
               12'b100100001011: data1 <=  20'h32641;
               12'b100100001100: data1 <=  20'h0f466;
               12'b100100001101: data1 <=  20'h6a707;
               12'b100100001110: data1 <=  20'h3c885;
               12'b100100001111: data1 <=  20'h22449;
               12'b100100010000: data1 <=  20'h3c885;
               12'b100100010001: data1 <=  20'h468a5;
               12'b100100010010: data1 <=  20'h54922;
               12'b100100010011: data1 <=  20'h06661;
               12'b100100010100: data1 <=  20'h72906;
               12'b100100010101: data1 <=  20'h4c908;
               12'b100100010110: data1 <=  20'h40542;
               12'b100100010111: data1 <=  20'h258c3;
               12'b100100011000: data1 <=  20'h73ce3;
               12'b100100011001: data1 <=  20'h714c3;
               12'b100100011010: data1 <=  20'h6d4c3;
               12'b100100011011: data1 <=  20'h775e4;
               12'b100100011100: data1 <=  20'h59cc8;
               12'b100100011101: data1 <=  20'h400e4;
               12'b100100011110: data1 <=  20'h3bcc3;
               12'b100100011111: data1 <=  20'h6b8c3;
               12'b100100100000: data1 <=  20'h35049;
               12'b100100100001: data1 <=  20'h27049;
               12'b100100100010: data1 <=  20'h3c866;
               12'b100100100011: data1 <=  20'h39466;
               12'b100100100100: data1 <=  20'h6dd22;
               12'b100100100101: data1 <=  20'h7d122;
               12'b100100100110: data1 <=  20'h80522;
               12'b100100100111: data1 <=  20'h7d922;
               12'b100100101000: data1 <=  20'h6be41;
               12'b100100101001: data1 <=  20'h6a641;
               12'b100100101010: data1 <=  20'h11c4b;
               12'b100100101011: data1 <=  20'h0cc4b;
               12'b100100101100: data1 <=  20'h03c38;
               12'b100100101101: data1 <=  20'h7fd04;
               12'b100100101110: data1 <=  20'h28c49;
               12'b100100101111: data1 <=  20'h3a0a7;
               12'b100100110000: data1 <=  20'h3bcc3;
               12'b100100110001: data1 <=  20'h390e3;
               12'b100100110010: data1 <=  20'h1e84a;
               12'b100100110011: data1 <=  20'h3a0c3;
               12'b100100110100: data1 <=  20'h030a7;
               12'b100100110101: data1 <=  20'h09126;
               12'b100100110110: data1 <=  20'h03c38;
               12'b100100110111: data1 <=  20'h02038;
               12'b100100111000: data1 <=  20'h4e467;
               12'b100100111001: data1 <=  20'h4d067;
               12'b100100111010: data1 <=  20'h218d3;
               12'b100100111011: data1 <=  20'h27866;
               12'b100100111100: data1 <=  20'h22466;
               12'b100100111101: data1 <=  20'h64ca4;
               12'b100100111110: data1 <=  20'h560a5;
               12'b100100111111: data1 <=  20'h514a5;
               12'b100101000000: data1 <=  20'h1e84a;
               12'b100101000001: data1 <=  20'h1904a;
               12'b100101000010: data1 <=  20'h2d8a4;
               12'b100101000011: data1 <=  20'h798e4;
               12'b100101000100: data1 <=  20'h474c3;
               12'b100101000101: data1 <=  20'h0cb01;
               12'b100101000110: data1 <=  20'h100ea;
               12'b100101000111: data1 <=  20'h51c49;
               12'b100101001000: data1 <=  20'h03453;
               12'b100101001001: data1 <=  20'h46ce3;
               12'b100101001010: data1 <=  20'h0a10a;
               12'b100101001011: data1 <=  20'h404e9;
               12'b100101001100: data1 <=  20'h798a5;
               12'b100101001101: data1 <=  20'h41466;
               12'b100101001110: data1 <=  20'h0a10a;
               12'b100101001111: data1 <=  20'h0690a;
               12'b100101010000: data1 <=  20'h42866;
               12'b100101010001: data1 <=  20'h3fc66;
               12'b100101010010: data1 <=  20'h288a4;
               12'b100101010011: data1 <=  20'h4c0c3;
               12'b100101010100: data1 <=  20'h2d582;
               12'b100101010101: data1 <=  20'h2e0a5;
               12'b100101010110: data1 <=  20'h10522;
               12'b100101010111: data1 <=  20'h20d65;
               12'b100101011000: data1 <=  20'h54486;
               12'b100101011001: data1 <=  20'h1ad22;
               12'b100101011010: data1 <=  20'h0e1a2;
               12'b100101011011: data1 <=  20'h28049;
               12'b100101011100: data1 <=  20'h35049;
               12'b100101011101: data1 <=  20'h7dd42;
               12'b100101011110: data1 <=  20'h5ee81;
               12'b100101011111: data1 <=  20'h6ad22;
               12'b100101100000: data1 <=  20'h03453;
               12'b100101100001: data1 <=  20'h02453;
               12'b100101100010: data1 <=  20'h1fac1;
               12'b100101100011: data1 <=  20'h0c922;
               12'b100101100100: data1 <=  20'h38709;
               12'b100101100101: data1 <=  20'h26604;
               12'b100101100110: data1 <=  20'h32e42;
               12'b100101100111: data1 <=  20'h0784a;
               12'b100101101000: data1 <=  20'h04066;
               12'b100101101001: data1 <=  20'h01466;
               12'b100101101010: data1 <=  20'h2e485;
               12'b100101101011: data1 <=  20'h20ce5;
               12'b100101101100: data1 <=  20'h0f942;
               12'b100101101101: data1 <=  20'h4ba61;
               12'b100101101110: data1 <=  20'h35049;
               12'b100101101111: data1 <=  20'h34849;
               12'b100101110000: data1 <=  20'h35449;
               12'b100101110001: data1 <=  20'h46469;
               12'b100101110010: data1 <=  20'h3a8c5;
               12'b100101110011: data1 <=  20'h5804a;
               12'b100101110100: data1 <=  20'h80903;
               12'b100101110101: data1 <=  20'h8a641;
               12'b100101110110: data1 <=  20'h1b8a6;
               12'b100101110111: data1 <=  20'h6ad82;
               12'b100101111000: data1 <=  20'h490c3;
               12'b100101111001: data1 <=  20'h4b942;
               12'b100101111010: data1 <=  20'h76f02;
               12'b100101111011: data1 <=  20'h72522;
               12'b100101111100: data1 <=  20'h0a84b;
               12'b100101111101: data1 <=  20'h0784b;
               12'b100101111110: data1 <=  20'h66d03;
               12'b100101111111: data1 <=  20'h08449;
               12'b100110000000: data1 <=  20'h41466;
               12'b100110000001: data1 <=  20'h334c3;
               12'b100110000010: data1 <=  20'h488a4;
               12'b100110000011: data1 <=  20'h45ca4;
               12'b100110000100: data1 <=  20'h29466;
               12'b100110000101: data1 <=  20'h27066;
               12'b100110000110: data1 <=  20'h3b4e4;
               12'b100110000111: data1 <=  20'h34467;
               12'b100110001000: data1 <=  20'h418c4;
               12'b100110001001: data1 <=  20'h20449;
               12'b100110001010: data1 <=  20'h4c206;
               12'b100110001011: data1 <=  20'h58cea;
               12'b100110001100: data1 <=  20'h5b106;
               12'b100110001101: data1 <=  20'h40c67;
               12'b100110001110: data1 <=  20'h22466;
               12'b100110001111: data1 <=  20'h1b832;
               12'b100110010000: data1 <=  20'h1c167;
               12'b100110010001: data1 <=  20'h32a41;
               12'b100110010010: data1 <=  20'h418c4;
               12'b100110010011: data1 <=  20'h21867;
               12'b100110010100: data1 <=  20'h54486;
               12'b100110010101: data1 <=  20'h53486;
               12'b100110010110: data1 <=  20'h5314b;
               12'b100110010111: data1 <=  20'h06834;
               12'b100110011000: data1 <=  20'h54922;
               12'b100110011001: data1 <=  20'h51d22;
               12'b100110011010: data1 <=  20'h6e122;
               12'b100110011011: data1 <=  20'h6a522;
               12'b100110011100: data1 <=  20'h03d2c;
               12'b100110011101: data1 <=  20'h400c4;
               12'b100110011110: data1 <=  20'h3a542;
               12'b100110011111: data1 <=  20'h38923;
               12'b100110100000: data1 <=  20'h2d641;
               12'b100110100001: data1 <=  20'h2e468;
               12'b100110100010: data1 <=  20'h4e04c;
               12'b100110100011: data1 <=  20'h5ea41;
               12'b100110100100: data1 <=  20'h6ec67;
               12'b100110100101: data1 <=  20'h57d42;
               12'b100110100110: data1 <=  20'h6ec67;
               12'b100110100111: data1 <=  20'h15833;
               12'b100110101000: data1 <=  20'h6ec67;
               12'b100110101001: data1 <=  20'h1a963;
               12'b100110101010: data1 <=  20'h6ec67;
               12'b100110101011: data1 <=  20'h33963;
               12'b100110101100: data1 <=  20'h2fc85;
               12'b100110101101: data1 <=  20'h1c153;
               12'b100110101110: data1 <=  20'h088e6;
               12'b100110101111: data1 <=  20'h20cc7;
               12'b100110110000: data1 <=  20'h02c49;
               12'b100110110001: data1 <=  20'h46485;
               12'b100110110010: data1 <=  20'h2fc85;
               12'b100110110011: data1 <=  20'h2cc85;
               12'b100110110100: data1 <=  20'h6ec67;
               12'b100110110101: data1 <=  20'h27885;
               12'b100110110110: data1 <=  20'h62469;
               12'b100110110111: data1 <=  20'h5e869;
               12'b100110111000: data1 <=  20'h42467;
               12'b100110111001: data1 <=  20'h40067;
               12'b100110111010: data1 <=  20'h624a4;
               12'b100110111011: data1 <=  20'h06466;
               12'b100110111100: data1 <=  20'h03466;
               12'b100110111101: data1 <=  20'h01ca6;
               12'b100110111110: data1 <=  20'h07508;
               12'b100110111111: data1 <=  20'h89a61;
               12'b100111000000: data1 <=  20'h3c122;
               12'b100111000001: data1 <=  20'h26522;
               12'b100111000010: data1 <=  20'h27cc5;
               12'b100111000011: data1 <=  20'h3a466;
               12'b100111000100: data1 <=  20'h1a5c3;
               12'b100111000101: data1 <=  20'h00c8a;
               12'b100111000110: data1 <=  20'h140e3;
               12'b100111000111: data1 <=  20'h28085;
               12'b100111001000: data1 <=  20'h0748e;
               12'b100111001001: data1 <=  20'h582c2;
               12'b100111001010: data1 <=  20'h7f0c3;
               12'b100111001011: data1 <=  20'h0ac67;
               12'b100111001100: data1 <=  20'h00c66;
               12'b100111001101: data1 <=  20'h4c226;
               12'b100111001110: data1 <=  20'h018c3;
               12'b100111001111: data1 <=  20'h2f122;
               12'b100111010000: data1 <=  20'h58942;
               12'b100111010001: data1 <=  20'h3b4a6;
               12'b100111010010: data1 <=  20'h08503;
               12'b100111010011: data1 <=  20'h48066;
               12'b100111010100: data1 <=  20'h46c66;
               12'b100111010101: data1 <=  20'h45a61;
               12'b100111010110: data1 <=  20'h1f4c3;
               12'b100111010111: data1 <=  20'h74142;
               12'b100111011000: data1 <=  20'h70942;
               12'b100111011001: data1 <=  20'h61522;
               12'b100111011010: data1 <=  20'h6a641;
               12'b100111011011: data1 <=  20'h6be41;
               12'b100111011100: data1 <=  20'h7d122;
               12'b100111011101: data1 <=  20'h61522;
               12'b100111011110: data1 <=  20'h0e849;
               12'b100111011111: data1 <=  20'h35c4c;
               12'b100111100000: data1 <=  20'h6c504;
               12'b100111100001: data1 <=  20'h7f8c3;
               12'b100111100010: data1 <=  20'h33c4c;
               12'b100111100011: data1 <=  20'h2d8c3;
               12'b100111100100: data1 <=  20'h28849;
               12'b100111100101: data1 <=  20'h7fcc3;
               12'b100111100110: data1 <=  20'h7ecc3;
               12'b100111100111: data1 <=  20'h0b86a;
               12'b100111101000: data1 <=  20'h0646a;
               12'b100111101001: data1 <=  20'h16849;
               12'b100111101010: data1 <=  20'h258c4;
               12'b100111101011: data1 <=  20'h3ccc3;
               12'b100111101100: data1 <=  20'h14849;
               12'b100111101101: data1 <=  20'h04049;
               12'b100111101110: data1 <=  20'h384c3;
               12'b100111101111: data1 <=  20'h1d88a;
               12'b100111110000: data1 <=  20'h1988a;
               12'b100111110001: data1 <=  20'h61522;
               12'b100111110010: data1 <=  20'h5e122;
               12'b100111110011: data1 <=  20'h600c3;
               12'b100111110100: data1 <=  20'h5f122;
               12'b100111110101: data1 <=  20'h07a41;
               12'b100111110110: data1 <=  20'h0f467;
               12'b100111110111: data1 <=  20'h09466;
               12'b100111111000: data1 <=  20'h08866;
               12'b100111111001: data1 <=  20'h288e3;
               12'b100111111010: data1 <=  20'h0f04d;
               12'b100111111011: data1 <=  20'h47cc3;
               12'b100111111100: data1 <=  20'h088cf;
               12'b100111111101: data1 <=  20'h03467;
               12'b100111111110: data1 <=  20'h26603;
               12'b100111111111: data1 <=  20'h2ec66;
               12'b101000000000: data1 <=  20'h2e049;
               12'b101000000001: data1 <=  20'h03458;
               12'b101000000010: data1 <=  20'h02458;
               12'b101000000011: data1 <=  20'h540a4;
               12'b101000000100: data1 <=  20'h6c122;
               12'b101000000101: data1 <=  20'h39a42;
               12'b101000000110: data1 <=  20'h534a4;
               12'b101000000111: data1 <=  20'h77e22;
               12'b101000001000: data1 <=  20'h12d27;
               12'b101000001001: data1 <=  20'h0cb01;
               12'b101000001010: data1 <=  20'h64241;
               12'b101000001011: data1 <=  20'h02c49;
               12'b101000001100: data1 <=  20'h391c6;
               12'b101000001101: data1 <=  20'h2ec66;
               12'b101000001110: data1 <=  20'h02849;
               12'b101000001111: data1 <=  20'h2884a;
               12'b101000010000: data1 <=  20'h01c49;
               12'b101000010001: data1 <=  20'h024e7;
               12'b101000010010: data1 <=  20'h47485;
               12'b101000010011: data1 <=  20'h2e868;
               12'b101000010100: data1 <=  20'h27c69;
               12'b101000010101: data1 <=  20'h5c485;
               12'b101000010110: data1 <=  20'h57c85;
               12'b101000010111: data1 <=  20'h03c85;
               12'b101000011000: data1 <=  20'h01485;
               12'b101000011001: data1 <=  20'h07cc5;
               12'b101000011010: data1 <=  20'h4d922;
               12'b101000011011: data1 <=  20'h35143;
               12'b101000011100: data1 <=  20'h28067;
               12'b101000011101: data1 <=  20'h22c88;
               12'b101000011110: data1 <=  20'h39104;
               12'b101000011111: data1 <=  20'h33ca4;
               12'b101000100000: data1 <=  20'h4cca4;
               12'b101000100001: data1 <=  20'h7a4a4;
               12'b101000100010: data1 <=  20'h01cc9;
               12'b101000100011: data1 <=  20'h1d8a4;
               12'b101000100100: data1 <=  20'h664c4;
               12'b101000100101: data1 <=  20'h2f0a6;
               12'b101000100110: data1 <=  20'h2d4a6;
               12'b101000100111: data1 <=  20'h280c7;
               12'b101000101000: data1 <=  20'h70a41;
               12'b101000101001: data1 <=  20'h71641;
               12'b101000101010: data1 <=  20'h1a04a;
               12'b101000101011: data1 <=  20'h04098;
               12'b101000101100: data1 <=  20'h0208f;
               12'b101000101101: data1 <=  20'h04098;
               12'b101000101110: data1 <=  20'h1acc9;
               12'b101000101111: data1 <=  20'h5b522;
               12'b101000110000: data1 <=  20'h39123;
               12'b101000110001: data1 <=  20'h368c3;
               12'b101000110010: data1 <=  20'h320c3;
               12'b101000110011: data1 <=  20'h2f122;
               12'b101000110100: data1 <=  20'h06cca;
               12'b101000110101: data1 <=  20'h04477;
               12'b101000110110: data1 <=  20'h5e049;
               12'b101000110111: data1 <=  20'h40942;
               12'b101000111000: data1 <=  20'h25943;
               12'b101000111001: data1 <=  20'h4ec85;
               12'b101000111010: data1 <=  20'h19433;
               12'b101000111011: data1 <=  20'h0b432;
               12'b101000111100: data1 <=  20'h07032;
               12'b101000111101: data1 <=  20'h40cc3;
               12'b101000111110: data1 <=  20'h1b4a9;
               12'b101000111111: data1 <=  20'h530e7;
               12'b101001000000: data1 <=  20'h53ce7;
               12'b101001000001: data1 <=  20'h60866;
               12'b101001000010: data1 <=  20'h58885;
               12'b101001000011: data1 <=  20'h79485;
               12'b101001000100: data1 <=  20'h64ca8;
               12'b101001000101: data1 <=  20'h4ed22;
               12'b101001000110: data1 <=  20'h4b122;
               12'b101001000111: data1 <=  20'h40183;
               12'b101001001000: data1 <=  20'h59ca4;
               12'b101001001001: data1 <=  20'h2ec66;
               12'b101001001010: data1 <=  20'h60449;
               12'b101001001011: data1 <=  20'h3c4e3;
               12'b101001001100: data1 <=  20'h08c56;
               12'b101001001101: data1 <=  20'h270e3;
               12'b101001001110: data1 <=  20'h76e61;
               12'b101001001111: data1 <=  20'h04478;
               12'b101001010000: data1 <=  20'h528a6;
               12'b101001010001: data1 <=  20'h290a7;
               12'b101001010010: data1 <=  20'h25c85;
               12'b101001010011: data1 <=  20'h274c5;
               12'b101001010100: data1 <=  20'h2e466;
               12'b101001010101: data1 <=  20'h358e7;
               12'b101001010110: data1 <=  20'h32ce7;
               12'b101001010111: data1 <=  20'h40da2;
               12'b101001011000: data1 <=  20'h0d466;
               12'b101001011001: data1 <=  20'h52e23;
               12'b101001011010: data1 <=  20'h51a23;
               12'b101001011011: data1 <=  20'h42903;
               12'b101001011100: data1 <=  20'h3e903;
               12'b101001011101: data1 <=  20'h3b585;
               12'b101001011110: data1 <=  20'h0e8a8;
               12'b101001011111: data1 <=  20'h0f0c8;
               12'b101001100000: data1 <=  20'h06522;
               12'b101001100001: data1 <=  20'h11c32;
               12'b101001100010: data1 <=  20'h13433;
               12'b101001100011: data1 <=  20'h37050;
               12'b101001100100: data1 <=  20'h32850;
               12'b101001100101: data1 <=  20'h7f162;
               12'b101001100110: data1 <=  20'h27885;
               12'b101001100111: data1 <=  20'h28485;
               12'b101001101000: data1 <=  20'h15066;
               12'b101001101001: data1 <=  20'h274c5;
               12'b101001101010: data1 <=  20'h35067;
               12'b101001101011: data1 <=  20'h0f466;
               12'b101001101100: data1 <=  20'h6c4c3;
               12'b101001101101: data1 <=  20'h0f466;
               12'b101001101110: data1 <=  20'h13d0a;
               12'b101001101111: data1 <=  20'h288a6;
               12'b101001110000: data1 <=  20'h258e4;
               12'b101001110001: data1 <=  20'h79d62;
               12'b101001110010: data1 <=  20'h2ccc4;
               12'b101001110011: data1 <=  20'h47c85;
               12'b101001110100: data1 <=  20'h09049;
               12'b101001110101: data1 <=  20'h03c36;
               12'b101001110110: data1 <=  20'h02036;
               12'b101001110111: data1 <=  20'h2f122;
               12'b101001111000: data1 <=  20'h2e485;
               12'b101001111001: data1 <=  20'h2ec66;
               12'b101001111010: data1 <=  20'h0252d;
               12'b101001111011: data1 <=  20'h04438;
               12'b101001111100: data1 <=  20'h01838;
               12'b101001111101: data1 <=  20'h794a4;
               12'b101001111110: data1 <=  20'h77641;
               12'b101001111111: data1 <=  20'h38e81;
               12'b101010000000: data1 <=  20'h33d22;
               12'b101010000001: data1 <=  20'h2ca65;
               12'b101010000010: data1 <=  20'h32a61;
               12'b101010000011: data1 <=  20'h35d22;
               12'b101010000100: data1 <=  20'h0e8c8;
               12'b101010000101: data1 <=  20'h3ace4;
               12'b101010000110: data1 <=  20'h1ac70;
               12'b101010000111: data1 <=  20'h36870;
               12'b101010001000: data1 <=  20'h32c70;
               12'b101010001001: data1 <=  20'h0504e;
               12'b101010001010: data1 <=  20'h0084e;
               12'b101010001011: data1 <=  20'h04456;
               12'b101010001100: data1 <=  20'h01456;
               12'b101010001101: data1 <=  20'h10894;
               12'b101010001110: data1 <=  20'h0d894;
               12'b101010001111: data1 <=  20'h28449;
               12'b101010010000: data1 <=  20'h03070;
               12'b101010010001: data1 <=  20'h2ec66;
               12'b101010010010: data1 <=  20'h19d23;
               12'b101010010011: data1 <=  20'h22904;
               12'b101010010100: data1 <=  20'h5dd42;
               12'b101010010101: data1 <=  20'h66122;
               12'b101010010110: data1 <=  20'h0ec66;
               12'b101010010111: data1 <=  20'h0b0a4;
               12'b101010011000: data1 <=  20'h2e066;
               12'b101010011001: data1 <=  20'h2d583;
               12'b101010011010: data1 <=  20'h21c86;
               12'b101010011011: data1 <=  20'h07885;
               12'b101010011100: data1 <=  20'h670c4;
               12'b101010011101: data1 <=  20'h58582;
               12'b101010011110: data1 <=  20'h744c3;
               12'b101010011111: data1 <=  20'h650c3;
               12'b101010100000: data1 <=  20'h4dce9;
               12'b101010100001: data1 <=  20'h3a8c3;
               12'b101010100010: data1 <=  20'h1a661;
               12'b101010100011: data1 <=  20'h0d8c3;
               12'b101010100100: data1 <=  20'h28449;
               12'b101010100101: data1 <=  20'h28049;
               12'b101010100110: data1 <=  20'h5b8a5;
               12'b101010100111: data1 <=  20'h584a5;
               12'b101010101000: data1 <=  20'h28ce3;
               12'b101010101001: data1 <=  20'h53467;
               12'b101010101010: data1 <=  20'h66105;
               12'b101010101011: data1 <=  20'h7f943;
               12'b101010101100: data1 <=  20'h46241;
               12'b101010101101: data1 <=  20'h2604a;
               12'b101010101110: data1 <=  20'h0d281;
               12'b101010101111: data1 <=  20'h5404b;
               12'b101010110000: data1 <=  20'h790c4;
               12'b101010110001: data1 <=  20'h600c3;
               12'b101010110010: data1 <=  20'h4c641;
               12'b101010110011: data1 <=  20'h329e2;
               12'b101010110100: data1 <=  20'h07e41;
               12'b101010110101: data1 <=  20'h01832;
               12'b101010110110: data1 <=  20'h17c4a;
               12'b101010110111: data1 <=  20'h1344a;
               12'b101010111000: data1 <=  20'h21c89;
               12'b101010111001: data1 <=  20'h21c89;
               12'b101010111010: data1 <=  20'h13a81;
               12'b101010111011: data1 <=  20'h1a5a2;
               12'b101010111100: data1 <=  20'h300e7;
               12'b101010111101: data1 <=  20'h2bce7;
               12'b101010111110: data1 <=  20'h470a6;
               12'b101010111111: data1 <=  20'h474a6;
               12'b101011000000: data1 <=  20'h4dc66;
               12'b101011000001: data1 <=  20'h6a641;
               12'b101011000010: data1 <=  20'h6be41;
               12'b101011000011: data1 <=  20'h45d25;
               12'b101011000100: data1 <=  20'h3a9e2;
               12'b101011000101: data1 <=  20'h26cc3;
               12'b101011000110: data1 <=  20'h1a983;
               12'b101011000111: data1 <=  20'h3a066;
               12'b101011001000: data1 <=  20'h2e9a2;
               12'b101011001001: data1 <=  20'h47d6d;
               12'b101011001010: data1 <=  20'h494c3;
               12'b101011001011: data1 <=  20'h44cc3;
               12'b101011001100: data1 <=  20'h2bf01;
               12'b101011001101: data1 <=  20'h2bd42;
               12'b101011001110: data1 <=  20'h33a41;
               12'b101011001111: data1 <=  20'h0c942;
               12'b101011010000: data1 <=  20'h05033;
               12'b101011010001: data1 <=  20'h268c8;
               12'b101011010010: data1 <=  20'h2ac49;
               12'b101011010011: data1 <=  20'h25c49;
               12'b101011010100: data1 <=  20'h8a641;
               12'b101011010101: data1 <=  20'h83522;
               12'b101011010110: data1 <=  20'h750c3;
               12'b101011010111: data1 <=  20'h7ed22;
               12'b101011011000: data1 <=  20'h684a4;
               12'b101011011001: data1 <=  20'h648a4;
               12'b101011011010: data1 <=  20'h04ca6;
               12'b101011011011: data1 <=  20'h000a6;
               12'b101011011100: data1 <=  20'h67d22;
               12'b101011011101: data1 <=  20'h64122;
               12'b101011011110: data1 <=  20'h67942;
               12'b101011011111: data1 <=  20'h64142;
               12'b101011100000: data1 <=  20'h78241;
               12'b101011100001: data1 <=  20'h76e41;
               12'b101011100010: data1 <=  20'h22526;
               12'b101011100011: data1 <=  20'h26ce3;
               12'b101011100100: data1 <=  20'h20665;
               12'b101011100101: data1 <=  20'h0d602;
               12'b101011100110: data1 <=  20'h4c10c;
               12'b101011100111: data1 <=  20'h154cf;
               12'b101011101000: data1 <=  20'h1d033;
               12'b101011101001: data1 <=  20'h1ac33;
               12'b101011101010: data1 <=  20'h5bc85;
               12'b101011101011: data1 <=  20'h58485;
               12'b101011101100: data1 <=  20'h4e066;
               12'b101011101101: data1 <=  20'h460c3;
               12'b101011101110: data1 <=  20'h22c85;
               12'b101011101111: data1 <=  20'h1a8c5;
               12'b101011110000: data1 <=  20'h35d25;
               12'b101011110001: data1 <=  20'h32125;
               12'b101011110010: data1 <=  20'h4e066;
               12'b101011110011: data1 <=  20'h5de41;
               12'b101011110100: data1 <=  20'h4e066;
               12'b101011110101: data1 <=  20'h4d466;
               12'b101011110110: data1 <=  20'h5f641;
               12'b101011110111: data1 <=  20'h25a41;
               12'b101011111000: data1 <=  20'h262c1;
               12'b101011111001: data1 <=  20'h01cea;
               12'b101011111010: data1 <=  20'h15cd1;
               12'b101011111011: data1 <=  20'h144d1;
               12'b101011111100: data1 <=  20'h4d10b;
               12'b101011111101: data1 <=  20'h52603;
               12'b101011111110: data1 <=  20'h4e0c4;
               12'b101011111111: data1 <=  20'h5a087;
               12'b101100000000: data1 <=  20'h43067;
               12'b101100000001: data1 <=  20'h3f467;
               12'b101100000010: data1 <=  20'h52e41;
               12'b101100000011: data1 <=  20'h3fd42;
               12'b101100000100: data1 <=  20'h54522;
               12'b101100000101: data1 <=  20'h51522;
               12'b101100000110: data1 <=  20'h0f832;
               12'b101100000111: data1 <=  20'h0f432;
               12'b101100001000: data1 <=  20'h4dc4a;
               12'b101100001001: data1 <=  20'h518c3;
               12'b101100001010: data1 <=  20'h3bd03;
               12'b101100001011: data1 <=  20'h3ed22;
               12'b101100001100: data1 <=  20'h3a202;
               12'b101100001101: data1 <=  20'h06641;
               12'b101100001110: data1 <=  20'h03049;
               12'b101100001111: data1 <=  20'h22466;
               12'b101100010000: data1 <=  20'h28849;
               12'b101100010001: data1 <=  20'h02849;
               12'b101100010010: data1 <=  20'h1b4c3;
               12'b101100010011: data1 <=  20'h13243;
               12'b101100010100: data1 <=  20'h19301;
               12'b101100010101: data1 <=  20'h65922;
               12'b101100010110: data1 <=  20'h3b485;
               12'b101100010111: data1 <=  20'h209a3;
               12'b101100011000: data1 <=  20'h2ce03;
               12'b101100011001: data1 <=  20'h2cdc3;
               12'b101100011010: data1 <=  20'h2dd22;
               12'b101100011011: data1 <=  20'h38a02;
               12'b101100011100: data1 <=  20'h349a3;
               12'b101100011101: data1 <=  20'h325a3;
               12'b101100011110: data1 <=  20'h1c183;
               12'b101100011111: data1 <=  20'h6a943;
               12'b101100100000: data1 <=  20'h71e41;
               12'b101100100001: data1 <=  20'h6a641;
               12'b101100100010: data1 <=  20'h79122;
               12'b101100100011: data1 <=  20'h7d562;
               12'b101100100100: data1 <=  20'h6c503;
               12'b101100100101: data1 <=  20'h46d05;
               12'b101100100110: data1 <=  20'h20a41;
               12'b101100100111: data1 <=  20'h344a5;
               12'b101100101000: data1 <=  20'h338c3;
               12'b101100101001: data1 <=  20'h26123;
               12'b101100101010: data1 <=  20'h28849;
               12'b101100101011: data1 <=  20'h21c66;
               12'b101100101100: data1 <=  20'h5b049;
               12'b101100101101: data1 <=  20'h59849;
               12'b101100101110: data1 <=  20'h0eca6;
               12'b101100101111: data1 <=  20'h0952c;
               12'b101100110000: data1 <=  20'h52a2b;
               12'b101100110001: data1 <=  20'h0d982;
               12'b101100110010: data1 <=  20'h3bd03;
               12'b101100110011: data1 <=  20'h3a8a9;
               12'b101100110100: data1 <=  20'h03849;
               12'b101100110101: data1 <=  20'h02049;
               12'b101100110110: data1 <=  20'h0904c;
               12'b101100110111: data1 <=  20'h461a2;
               12'b101100111000: data1 <=  20'h39a61;
               12'b101100111001: data1 <=  20'h538c4;
               12'b101100111010: data1 <=  20'h5a485;
               12'b101100111011: data1 <=  20'h00867;
               12'b101100111100: data1 <=  20'h0ac67;
               12'b101100111101: data1 <=  20'h07067;
               12'b101100111110: data1 <=  20'h80122;
               12'b101100111111: data1 <=  20'h0144a;
               12'b101101000000: data1 <=  20'h37086;
               12'b101101000001: data1 <=  20'h32086;
               12'b101101000010: data1 <=  20'h55ca4;
               12'b101101000011: data1 <=  20'h518a4;
               12'b101101000100: data1 <=  20'h55085;
               12'b101101000101: data1 <=  20'h52885;
               12'b101101000110: data1 <=  20'h5f604;
               12'b101101000111: data1 <=  20'h5e604;
               12'b101101001000: data1 <=  20'h614e3;
               12'b101101001001: data1 <=  20'h34867;
               12'b101101001010: data1 <=  20'h54922;
               12'b101101001011: data1 <=  20'h52223;
               12'b101101001100: data1 <=  20'h54905;
               12'b101101001101: data1 <=  20'h52105;
               12'b101101001110: data1 <=  20'h5b8a4;
               12'b101101001111: data1 <=  20'h70963;
               12'b101101010000: data1 <=  20'h64184;
               12'b101101010001: data1 <=  20'h800c3;
               12'b101101010010: data1 <=  20'h50466;
               12'b101101010011: data1 <=  20'h4b066;
               12'b101101010100: data1 <=  20'h7a922;
               12'b101101010101: data1 <=  20'h25d65;
               12'b101101010110: data1 <=  20'h7a922;
               12'b101101010111: data1 <=  20'h76e41;
               12'b101101011000: data1 <=  20'h64e61;
               12'b101101011001: data1 <=  20'h57a41;
               12'b101101011010: data1 <=  20'h7a922;
               12'b101101011011: data1 <=  20'h76d22;
               12'b101101011100: data1 <=  20'h79d22;
               12'b101101011101: data1 <=  20'h77922;
               12'b101101011110: data1 <=  20'h10c34;
               12'b101101011111: data1 <=  20'h6a704;
               12'b101101100000: data1 <=  20'h0946b;
               default: data1 <= 0;
           endcase
        end

endmodule: rect1_rom
