module sqrt_rom_mem
  #(
     W_DATA = 16,
     DEPTH = 64,
     W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input ena,
     input [W_ADDR-1:0] addra,
     output [W_DATA-1:0] doa

     );

     logic [W_DATA-1:0] mem [DEPTH-1:0];

     always_ff @(posedge clk)
        begin
           if(ena)
              doa = mem[addra];
        end

     initial begin
         mem[0] = 16'h0000;
         mem[1] = 16'h0b50;
         mem[2] = 16'h1000;
         mem[3] = 16'h1398;
         mem[4] = 16'h16a0;
         mem[5] = 16'h194c;
         mem[6] = 16'h1bb6;
         mem[7] = 16'h1dee;
         mem[8] = 16'h2000;
         mem[9] = 16'h21f0;
         mem[10] = 16'h23c6;
         mem[11] = 16'h2585;
         mem[12] = 16'h2731;
         mem[13] = 16'h28ca;
         mem[14] = 16'h2a54;
         mem[15] = 16'h2bd1;
         mem[16] = 16'h2d41;
         mem[17] = 16'h2ea5;
         mem[18] = 16'h3000;
         mem[19] = 16'h3150;
         mem[20] = 16'h3298;
         mem[21] = 16'h33d8;
         mem[22] = 16'h3510;
         mem[23] = 16'h3642;
         mem[24] = 16'h376c;
         mem[25] = 16'h3891;
         mem[26] = 16'h39b0;
         mem[27] = 16'h3ac9;
         mem[28] = 16'h3bdd;
         mem[29] = 16'h3ced;
         mem[30] = 16'h3df7;
         mem[31] = 16'h3efd;
         mem[32] = 16'h4000;
         mem[33] = 16'h40fe;
         mem[34] = 16'h41f8;
         mem[35] = 16'h42ee;
         mem[36] = 16'h43e1;
         mem[37] = 16'h44d1;
         mem[38] = 16'h45be;
         mem[39] = 16'h46a7;
         mem[40] = 16'h478d;
         mem[41] = 16'h4871;
         mem[42] = 16'h4952;
         mem[43] = 16'h4a30;
         mem[44] = 16'h4b0b;
         mem[45] = 16'h4be5;
         mem[46] = 16'h4cbb;
         mem[47] = 16'h4d90;
         mem[48] = 16'h4e62;
         mem[49] = 16'h4f32;
         mem[50] = 16'h5000;
         mem[51] = 16'h50cb;
         mem[52] = 16'h5195;
         mem[53] = 16'h525d;
         mem[54] = 16'h5323;
         mem[55] = 16'h53e7;
         mem[56] = 16'h54a9;
         mem[57] = 16'h556a;
         mem[58] = 16'h5629;
         mem[59] = 16'h56e6;
         mem[60] = 16'h57a2;
         mem[61] = 16'h585c;
         mem[62] = 16'h5915;
         mem[63] = 16'h59cc;
         mem[64] = 16'h5a82;
         mem[65] = 16'h5b36;
         mem[66] = 16'h5be9;
         mem[67] = 16'h5c9b;
         mem[68] = 16'h5d4b;
         mem[69] = 16'h5dfa;
         mem[70] = 16'h5ea8;
         mem[71] = 16'h5f54;
         mem[72] = 16'h6000;
         mem[73] = 16'h60aa;
         mem[74] = 16'h6152;
         mem[75] = 16'h61fa;
         mem[76] = 16'h62a1;
         mem[77] = 16'h6347;
         mem[78] = 16'h63eb;
         mem[79] = 16'h648e;
         mem[80] = 16'h6531;
         mem[81] = 16'h65d2;
         mem[82] = 16'h6673;
         mem[83] = 16'h6712;
         mem[84] = 16'h67b1;
         mem[85] = 16'h684e;
         mem[86] = 16'h68eb;
         mem[87] = 16'h6986;
         mem[88] = 16'h6a21;
         mem[89] = 16'h6abb;
         mem[90] = 16'h6b54;
         mem[91] = 16'h6bed;
         mem[92] = 16'h6c84;
         mem[93] = 16'h6d1a;
         mem[94] = 16'h6db0;
         mem[95] = 16'h6e45;
         mem[96] = 16'h6ed9;
         mem[97] = 16'h6f6d;
         mem[98] = 16'h7000;
         mem[99] = 16'h7091;
         mem[100] = 16'h7123;
         mem[101] = 16'h71b3;
         mem[102] = 16'h7243;
         mem[103] = 16'h72d2;
         mem[104] = 16'h7360;
         mem[105] = 16'h73ee;
         mem[106] = 16'h747b;
         mem[107] = 16'h7507;
         mem[108] = 16'h7593;
         mem[109] = 16'h761e;
         mem[110] = 16'h76a8;
         mem[111] = 16'h7732;
         mem[112] = 16'h77bb;
         mem[113] = 16'h7844;
         mem[114] = 16'h78cc;
         mem[115] = 16'h7953;
         mem[116] = 16'h79da;
         mem[117] = 16'h7a60;
         mem[118] = 16'h7ae5;
         mem[119] = 16'h7b6b;
         mem[120] = 16'h7bef;
         mem[121] = 16'h7c73;
         mem[122] = 16'h7cf6;
         mem[123] = 16'h7d79;
         mem[124] = 16'h7dfb;
         mem[125] = 16'h7e7d;
         mem[126] = 16'h7efe;
         mem[127] = 16'h7f7f;
         mem[128] = 16'h8000;
         mem[129] = 16'h807f;
         mem[130] = 16'h80ff;
         mem[131] = 16'h817d;
         mem[132] = 16'h81fc;
         mem[133] = 16'h8279;
         mem[134] = 16'h82f7;
         mem[135] = 16'h8374;
         mem[136] = 16'h83f0;
         mem[137] = 16'h846c;
         mem[138] = 16'h84e7;
         mem[139] = 16'h8562;
         mem[140] = 16'h85dd;
         mem[141] = 16'h8657;
         mem[142] = 16'h86d1;
         mem[143] = 16'h874a;
         mem[144] = 16'h87c3;
         mem[145] = 16'h883c;
         mem[146] = 16'h88b4;
         mem[147] = 16'h892b;
         mem[148] = 16'h89a3;
         mem[149] = 16'h8a19;
         mem[150] = 16'h8a90;
         mem[151] = 16'h8b06;
         mem[152] = 16'h8b7c;
         mem[153] = 16'h8bf1;
         mem[154] = 16'h8c66;
         mem[155] = 16'h8cda;
         mem[156] = 16'h8d4e;
         mem[157] = 16'h8dc2;
         mem[158] = 16'h8e36;
         mem[159] = 16'h8ea9;
         mem[160] = 16'h8f1b;
         mem[161] = 16'h8f8e;
         mem[162] = 16'h9000;
         mem[163] = 16'h9071;
         mem[164] = 16'h90e2;
         mem[165] = 16'h9153;
         mem[166] = 16'h91c4;
         mem[167] = 16'h9234;
         mem[168] = 16'h92a4;
         mem[169] = 16'h9314;
         mem[170] = 16'h9383;
         mem[171] = 16'h93f2;
         mem[172] = 16'h9460;
         mem[173] = 16'h94cf;
         mem[174] = 16'h953c;
         mem[175] = 16'h95aa;
         mem[176] = 16'h9617;
         mem[177] = 16'h9684;
         mem[178] = 16'h96f1;
         mem[179] = 16'h975d;
         mem[180] = 16'h97ca;
         mem[181] = 16'h9835;
         mem[182] = 16'h98a1;
         mem[183] = 16'h990c;
         mem[184] = 16'h9977;
         mem[185] = 16'h99e2;
         mem[186] = 16'h9a4c;
         mem[187] = 16'h9ab6;
         mem[188] = 16'h9b20;
         mem[189] = 16'h9b89;
         mem[190] = 16'h9bf2;
         mem[191] = 16'h9c5b;
         mem[192] = 16'h9cc4;
         mem[193] = 16'h9d2c;
         mem[194] = 16'h9d94;
         mem[195] = 16'h9dfc;
         mem[196] = 16'h9e64;
         mem[197] = 16'h9ecb;
         mem[198] = 16'h9f32;
         mem[199] = 16'h9f99;
         mem[200] = 16'ha000;
         mem[201] = 16'ha066;
         mem[202] = 16'ha0cc;
         mem[203] = 16'ha132;
         mem[204] = 16'ha197;
         mem[205] = 16'ha1fc;
         mem[206] = 16'ha261;
         mem[207] = 16'ha2c6;
         mem[208] = 16'ha32b;
         mem[209] = 16'ha38f;
         mem[210] = 16'ha3f3;
         mem[211] = 16'ha457;
         mem[212] = 16'ha4ba;
         mem[213] = 16'ha51e;
         mem[214] = 16'ha581;
         mem[215] = 16'ha5e4;
         mem[216] = 16'ha646;
         mem[217] = 16'ha6a9;
         mem[218] = 16'ha70b;
         mem[219] = 16'ha76d;
         mem[220] = 16'ha7cf;
         mem[221] = 16'ha830;
         mem[222] = 16'ha892;
         mem[223] = 16'ha8f3;
         mem[224] = 16'ha953;
         mem[225] = 16'ha9b4;
         mem[226] = 16'haa15;
         mem[227] = 16'haa75;
         mem[228] = 16'haad5;
         mem[229] = 16'hab35;
         mem[230] = 16'hab94;
         mem[231] = 16'habf4;
         mem[232] = 16'hac53;
         mem[233] = 16'hacb2;
         mem[234] = 16'had11;
         mem[235] = 16'had6f;
         mem[236] = 16'hadcd;
         mem[237] = 16'hae2c;
         mem[238] = 16'hae8a;
         mem[239] = 16'haee7;
         mem[240] = 16'haf45;
         mem[241] = 16'hafa2;
         mem[242] = 16'hb000;
         mem[243] = 16'hb05c;
         mem[244] = 16'hb0b9;
         mem[245] = 16'hb116;
         mem[246] = 16'hb172;
         mem[247] = 16'hb1cf;
         mem[248] = 16'hb22b;
         mem[249] = 16'hb286;
         mem[250] = 16'hb2e2;
         mem[251] = 16'hb33e;
         mem[252] = 16'hb399;
         mem[253] = 16'hb3f4;
         mem[254] = 16'hb44f;
         mem[255] = 16'hb4aa;
     end


endmodule: sqrt_rom_mem
