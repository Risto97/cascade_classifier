module rect0_rom
  #(
     parameter W_DATA = 20,
     parameter W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );
     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               12'b000000000000: data1 <=  20'h1a989;
               12'b000000000001: data1 <=  20'h1a987;
               12'b000000000010: data1 <=  20'h39249;
               12'b000000000011: data1 <=  20'h72926;
               12'b000000000100: data1 <=  20'h20093;
               12'b000000000101: data1 <=  20'h20d90;
               12'b000000000110: data1 <=  20'h33586;
               12'b000000000111: data1 <=  20'h5a48a;
               12'b000000001000: data1 <=  20'h010e6;
               12'b000000001001: data1 <=  20'h27186;
               12'b000000001010: data1 <=  20'h1a987;
               12'b000000001011: data1 <=  20'h3266c;
               12'b000000001100: data1 <=  20'h0cb03;
               12'b000000001101: data1 <=  20'h3a8cf;
               12'b000000001110: data1 <=  20'h26dca;
               12'b000000001111: data1 <=  20'h015c9;
               12'b000000010000: data1 <=  20'h48126;
               12'b000000010001: data1 <=  20'h210ca;
               12'b000000010010: data1 <=  20'h348ca;
               12'b000000010011: data1 <=  20'h1fc89;
               12'b000000010100: data1 <=  20'h048cb;
               12'b000000010101: data1 <=  20'h25b0d;
               12'b000000010110: data1 <=  20'h27cc9;
               12'b000000010111: data1 <=  20'h72546;
               12'b000000011000: data1 <=  20'h2d1cc;
               12'b000000011001: data1 <=  20'h12f03;
               12'b000000011010: data1 <=  20'h335e6;
               12'b000000011011: data1 <=  20'h27cae;
               12'b000000011100: data1 <=  20'h218ca;
               12'b000000011101: data1 <=  20'h2706c;
               12'b000000011110: data1 <=  20'h84243;
               12'b000000011111: data1 <=  20'h26da6;
               12'b000000100000: data1 <=  20'h0accf;
               12'b000000100001: data1 <=  20'h068cf;
               12'b000000100010: data1 <=  20'h3230f;
               12'b000000100011: data1 <=  20'h26dcc;
               12'b000000100100: data1 <=  20'h4baac;
               12'b000000100101: data1 <=  20'h0848a;
               12'b000000100110: data1 <=  20'h51e8a;
               12'b000000100111: data1 <=  20'h064cd;
               12'b000000101000: data1 <=  20'h1188d;
               12'b000000101001: data1 <=  20'h1f6d3;
               12'b000000101010: data1 <=  20'h1d8c9;
               12'b000000101011: data1 <=  20'h12ccb;
               12'b000000101100: data1 <=  20'h09489;
               12'b000000101101: data1 <=  20'h25a63;
               12'b000000101110: data1 <=  20'h09489;
               12'b000000101111: data1 <=  20'h08489;
               12'b000000110000: data1 <=  20'h209ce;
               12'b000000110001: data1 <=  20'h3ee42;
               12'b000000110010: data1 <=  20'h5588b;
               12'b000000110011: data1 <=  20'h190c9;
               12'b000000110100: data1 <=  20'h1a989;
               12'b000000110101: data1 <=  20'h20d86;
               12'b000000110110: data1 <=  20'h06705;
               12'b000000110111: data1 <=  20'h3fa46;
               12'b000000111000: data1 <=  20'h6ad86;
               12'b000000111001: data1 <=  20'h1788d;
               12'b000000111010: data1 <=  20'h1308d;
               12'b000000111011: data1 <=  20'h06717;
               12'b000000111100: data1 <=  20'h2c10c;
               12'b000000111101: data1 <=  20'h2f46e;
               12'b000000111110: data1 <=  20'h4be06;
               12'b000000111111: data1 <=  20'h27186;
               12'b000001000000: data1 <=  20'h2dccc;
               12'b000001000001: data1 <=  20'h61926;
               12'b000001000010: data1 <=  20'h6aa43;
               12'b000001000011: data1 <=  20'h1a20c;
               12'b000001000100: data1 <=  20'h06494;
               12'b000001000101: data1 <=  20'h00e42;
               12'b000001000110: data1 <=  20'h1fa8e;
               12'b000001000111: data1 <=  20'h335cc;
               12'b000001001000: data1 <=  20'h584e9;
               12'b000001001001: data1 <=  20'h61526;
               12'b000001001010: data1 <=  20'h5e126;
               12'b000001001011: data1 <=  20'h2850a;
               12'b000001001100: data1 <=  20'h209ce;
               12'b000001001101: data1 <=  20'h01985;
               12'b000001001110: data1 <=  20'h024c9;
               12'b000001001111: data1 <=  20'h27cc9;
               12'b000001010000: data1 <=  20'h01cc9;
               12'b000001010001: data1 <=  20'h280c9;
               12'b000001010010: data1 <=  20'h278c9;
               12'b000001010011: data1 <=  20'h32e44;
               12'b000001010100: data1 <=  20'h01989;
               12'b000001010101: data1 <=  20'h00306;
               12'b000001010110: data1 <=  20'h2ce0c;
               12'b000001010111: data1 <=  20'h284c6;
               12'b000001011000: data1 <=  20'h7d303;
               12'b000001011001: data1 <=  20'h28489;
               12'b000001011010: data1 <=  20'h525e4;
               12'b000001011011: data1 <=  20'h28489;
               12'b000001011100: data1 <=  20'h27c89;
               12'b000001011101: data1 <=  20'h4d4cc;
               12'b000001011110: data1 <=  20'h89e42;
               12'b000001011111: data1 <=  20'h2e48a;
               12'b000001100000: data1 <=  20'h2d50a;
               12'b000001100001: data1 <=  20'h27546;
               12'b000001100010: data1 <=  20'h57944;
               12'b000001100011: data1 <=  20'h72242;
               12'b000001100100: data1 <=  20'h06ac3;
               12'b000001100101: data1 <=  20'h65a43;
               12'b000001100110: data1 <=  20'h198cf;
               12'b000001100111: data1 <=  20'h1e08a;
               12'b000001101000: data1 <=  20'h1908a;
               12'b000001101001: data1 <=  20'h64a86;
               12'b000001101010: data1 <=  20'h4b109;
               12'b000001101011: data1 <=  20'h030c9;
               12'b000001101100: data1 <=  20'h3fcc6;
               12'b000001101101: data1 <=  20'h34d86;
               12'b000001101110: data1 <=  20'h32186;
               12'b000001101111: data1 <=  20'h030c9;
               12'b000001110000: data1 <=  20'h018c9;
               12'b000001110001: data1 <=  20'h59926;
               12'b000001110010: data1 <=  20'h64126;
               12'b000001110011: data1 <=  20'h348ca;
               12'b000001110100: data1 <=  20'h77983;
               12'b000001110101: data1 <=  20'h3f282;
               12'b000001110110: data1 <=  20'h38e4c;
               12'b000001110111: data1 <=  20'h00e58;
               12'b000001111000: data1 <=  20'h26dca;
               12'b000001111001: data1 <=  20'h2194c;
               12'b000001111010: data1 <=  20'h2058c;
               12'b000001111011: data1 <=  20'h58a43;
               12'b000001111100: data1 <=  20'h52d08;
               12'b000001111101: data1 <=  20'h64e46;
               12'b000001111110: data1 <=  20'h000c6;
               12'b000001111111: data1 <=  20'h27192;
               12'b000010000000: data1 <=  20'h07c8e;
               12'b000010000001: data1 <=  20'h0d662;
               12'b000010000010: data1 <=  20'h326cd;
               12'b000010000011: data1 <=  20'h3a564;
               12'b000010000100: data1 <=  20'h4b1ea;
               12'b000010000101: data1 <=  20'h67186;
               12'b000010000110: data1 <=  20'h64186;
               12'b000010000111: data1 <=  20'h0b0ac;
               12'b000010001000: data1 <=  20'h0cb04;
               12'b000010001001: data1 <=  20'h33984;
               12'b000010001010: data1 <=  20'h21126;
               12'b000010001011: data1 <=  20'h6c8c6;
               12'b000010001100: data1 <=  20'h2becf;
               12'b000010001101: data1 <=  20'h07629;
               12'b000010001110: data1 <=  20'h210ca;
               12'b000010001111: data1 <=  20'h0acc8;
               12'b000010010000: data1 <=  20'h064c7;
               12'b000010010001: data1 <=  20'h048d6;
               12'b000010010010: data1 <=  20'h000d6;
               12'b000010010011: data1 <=  20'h2fd10;
               12'b000010010100: data1 <=  20'h3f266;
               12'b000010010101: data1 <=  20'h3a8cc;
               12'b000010010110: data1 <=  20'h5e626;
               12'b000010010111: data1 <=  20'h2f46e;
               12'b000010011000: data1 <=  20'h26d0a;
               12'b000010011001: data1 <=  20'h35d2b;
               12'b000010011010: data1 <=  20'h3212b;
               12'b000010011011: data1 <=  20'h27952;
               12'b000010011100: data1 <=  20'h2d86e;
               12'b000010011101: data1 <=  20'h57b08;
               12'b000010011110: data1 <=  20'h3ee4e;
               12'b000010011111: data1 <=  20'h4e8c6;
               12'b000010100000: data1 <=  20'h01d50;
               12'b000010100001: data1 <=  20'h02926;
               12'b000010100010: data1 <=  20'h13e04;
               12'b000010100011: data1 <=  20'h02926;
               12'b000010100100: data1 <=  20'h06a84;
               12'b000010100101: data1 <=  20'h02926;
               12'b000010100110: data1 <=  20'h01526;
               12'b000010100111: data1 <=  20'h72946;
               12'b000010101000: data1 <=  20'h144c9;
               12'b000010101001: data1 <=  20'h14986;
               12'b000010101010: data1 <=  20'h3ea43;
               12'b000010101011: data1 <=  20'h3eec3;
               12'b000010101100: data1 <=  20'h46108;
               12'b000010101101: data1 <=  20'h47cc6;
               12'b000010101110: data1 <=  20'h464c6;
               12'b000010101111: data1 <=  20'h40566;
               12'b000010110000: data1 <=  20'h51704;
               12'b000010110001: data1 <=  20'h19acc;
               12'b000010110010: data1 <=  20'h00a91;
               12'b000010110011: data1 <=  20'h03858;
               12'b000010110100: data1 <=  20'h02058;
               12'b000010110101: data1 <=  20'h09c56;
               12'b000010110110: data1 <=  20'h08456;
               12'b000010110111: data1 <=  20'h29c72;
               12'b000010111000: data1 <=  20'h59126;
               12'b000010111001: data1 <=  20'h5ad24;
               12'b000010111010: data1 <=  20'h71643;
               12'b000010111011: data1 <=  20'h1b512;
               12'b000010111100: data1 <=  20'h6a643;
               12'b000010111101: data1 <=  20'h0c984;
               12'b000010111110: data1 <=  20'h339c6;
               12'b000010111111: data1 <=  20'h210c6;
               12'b000011000000: data1 <=  20'h21cd0;
               12'b000011000001: data1 <=  20'h19530;
               12'b000011000010: data1 <=  20'h01649;
               12'b000011000011: data1 <=  20'h600a8;
               12'b000011000100: data1 <=  20'h05089;
               12'b000011000101: data1 <=  20'h00a43;
               12'b000011000110: data1 <=  20'h8ae62;
               12'b000011000111: data1 <=  20'h00089;
               12'b000011001000: data1 <=  20'h26e72;
               12'b000011001001: data1 <=  20'h064c9;
               12'b000011001010: data1 <=  20'h20dcc;
               12'b000011001011: data1 <=  20'h06682;
               12'b000011001100: data1 <=  20'h0cec3;
               12'b000011001101: data1 <=  20'h328e9;
               12'b000011001110: data1 <=  20'h4bac4;
               12'b000011001111: data1 <=  20'h4b2c4;
               12'b000011010000: data1 <=  20'h2e0cb;
               12'b000011010001: data1 <=  20'h08126;
               12'b000011010010: data1 <=  20'h0f48a;
               12'b000011010011: data1 <=  20'h1a98c;
               12'b000011010100: data1 <=  20'h0accf;
               12'b000011010101: data1 <=  20'h5ea43;
               12'b000011010110: data1 <=  20'h23cc9;
               12'b000011010111: data1 <=  20'h1fa06;
               12'b000011011000: data1 <=  20'h02cc9;
               12'b000011011001: data1 <=  20'h1930e;
               12'b000011011010: data1 <=  20'h0348d;
               12'b000011011011: data1 <=  20'h01c8d;
               12'b000011011100: data1 <=  20'h284c9;
               12'b000011011101: data1 <=  20'h2dcc9;
               12'b000011011110: data1 <=  20'h6d926;
               12'b000011011111: data1 <=  20'h711c6;
               12'b000011100000: data1 <=  20'h71644;
               12'b000011100001: data1 <=  20'h7d1e4;
               12'b000011100010: data1 <=  20'h601e9;
               12'b000011100011: data1 <=  20'h1a204;
               12'b000011100100: data1 <=  20'h27546;
               12'b000011100101: data1 <=  20'h579ea;
               12'b000011100110: data1 <=  20'h3a14e;
               12'b000011100111: data1 <=  20'h274c9;
               12'b000011101000: data1 <=  20'h26643;
               12'b000011101001: data1 <=  20'h3ea43;
               12'b000011101010: data1 <=  20'h64e44;
               12'b000011101011: data1 <=  20'h269c6;
               12'b000011101100: data1 <=  20'h03452;
               12'b000011101101: data1 <=  20'h02452;
               12'b000011101110: data1 <=  20'h2d1ea;
               12'b000011101111: data1 <=  20'h7d6a4;
               12'b000011110000: data1 <=  20'h21cb2;
               12'b000011110001: data1 <=  20'h0cb06;
               12'b000011110010: data1 <=  20'h06ac8;
               12'b000011110011: data1 <=  20'h011e9;
               12'b000011110100: data1 <=  20'h00313;
               12'b000011110101: data1 <=  20'h83e43;
               12'b000011110110: data1 <=  20'h2e144;
               12'b000011110111: data1 <=  20'h2d144;
               12'b000011111000: data1 <=  20'h364d0;
               12'b000011111001: data1 <=  20'h5e284;
               12'b000011111010: data1 <=  20'h61546;
               12'b000011111011: data1 <=  20'h00e09;
               12'b000011111100: data1 <=  20'h294ef;
               12'b000011111101: data1 <=  20'h088cd;
               12'b000011111110: data1 <=  20'h10cce;
               12'b000011111111: data1 <=  20'h5858a;
               12'b000100000000: data1 <=  20'h27546;
               12'b000100000001: data1 <=  20'h0ccce;
               12'b000100000010: data1 <=  20'h1b8ac;
               12'b000100000011: data1 <=  20'h6a705;
               12'b000100000100: data1 <=  20'h2f8ac;
               12'b000100000101: data1 <=  20'h070cc;
               12'b000100000110: data1 <=  20'h544c6;
               12'b000100000111: data1 <=  20'h52cc6;
               12'b000100001000: data1 <=  20'h29070;
               12'b000100001001: data1 <=  20'h4b5a6;
               12'b000100001010: data1 <=  20'h09889;
               12'b000100001011: data1 <=  20'h01d26;
               12'b000100001100: data1 <=  20'h0f8c9;
               12'b000100001101: data1 <=  20'h0e0c9;
               12'b000100001110: data1 <=  20'h72186;
               12'b000100001111: data1 <=  20'h274c9;
               12'b000100010000: data1 <=  20'h2d983;
               12'b000100010001: data1 <=  20'h14d15;
               12'b000100010010: data1 <=  20'h1ad4c;
               12'b000100010011: data1 <=  20'h064c9;
               12'b000100010100: data1 <=  20'h10454;
               12'b000100010101: data1 <=  20'h12cc9;
               12'b000100010110: data1 <=  20'h16855;
               12'b000100010111: data1 <=  20'h01c57;
               12'b000100011000: data1 <=  20'h35d24;
               12'b000100011001: data1 <=  20'h32124;
               12'b000100011010: data1 <=  20'h59926;
               12'b000100011011: data1 <=  20'h57926;
               12'b000100011100: data1 <=  20'h3f644;
               12'b000100011101: data1 <=  20'h00313;
               12'b000100011110: data1 <=  20'h0890c;
               12'b000100011111: data1 <=  20'h2808a;
               12'b000100100000: data1 <=  20'h3a14c;
               12'b000100100001: data1 <=  20'h01473;
               12'b000100100010: data1 <=  20'h038ca;
               12'b000100100011: data1 <=  20'h008cc;
               12'b000100100100: data1 <=  20'h44f02;
               12'b000100100101: data1 <=  20'h395a4;
               12'b000100100110: data1 <=  20'h344c9;
               12'b000100100111: data1 <=  20'h4b204;
               12'b000100101000: data1 <=  20'h4f8c9;
               12'b000100101001: data1 <=  20'h4b0c9;
               12'b000100101010: data1 <=  20'h2dd44;
               12'b000100101011: data1 <=  20'h2dcc9;
               12'b000100101100: data1 <=  20'h02cc9;
               12'b000100101101: data1 <=  20'h01cc9;
               12'b000100101110: data1 <=  20'h15ccf;
               12'b000100101111: data1 <=  20'h144cf;
               12'b000100110000: data1 <=  20'h10524;
               12'b000100110001: data1 <=  20'h3fcc7;
               12'b000100110010: data1 <=  20'h59cca;
               12'b000100110011: data1 <=  20'h530a8;
               12'b000100110100: data1 <=  20'h22c70;
               12'b000100110101: data1 <=  20'h6ae43;
               12'b000100110110: data1 <=  20'h71e63;
               12'b000100110111: data1 <=  20'h024c9;
               12'b000100111000: data1 <=  20'h1c072;
               12'b000100111001: data1 <=  20'h1b472;
               12'b000100111010: data1 <=  20'h13a49;
               12'b000100111011: data1 <=  20'h07cce;
               12'b000100111100: data1 <=  20'h67126;
               12'b000100111101: data1 <=  20'h13290;
               12'b000100111110: data1 <=  20'h224cc;
               12'b000100111111: data1 <=  20'h0ced0;
               12'b000101000000: data1 <=  20'h5a0aa;
               12'b000101000001: data1 <=  20'h84243;
               12'b000101000010: data1 <=  20'h5a0ca;
               12'b000101000011: data1 <=  20'h0cb04;
               12'b000101000100: data1 <=  20'h1a989;
               12'b000101000101: data1 <=  20'h27185;
               12'b000101000110: data1 <=  20'h335cc;
               12'b000101000111: data1 <=  20'h5890a;
               12'b000101001000: data1 <=  20'h284ae;
               12'b000101001001: data1 <=  20'h27470;
               12'b000101001010: data1 <=  20'h2ca48;
               12'b000101001011: data1 <=  20'h13682;
               12'b000101001100: data1 <=  20'h4be66;
               12'b000101001101: data1 <=  20'h278c9;
               12'b000101001110: data1 <=  20'h298ce;
               12'b000101001111: data1 <=  20'h3a0cc;
               12'b000101010000: data1 <=  20'h2a0d2;
               12'b000101010001: data1 <=  20'h258d2;
               12'b000101010010: data1 <=  20'h110c9;
               12'b000101010011: data1 <=  20'h715e6;
               12'b000101010100: data1 <=  20'h110c9;
               12'b000101010101: data1 <=  20'h0c8c9;
               12'b000101010110: data1 <=  20'h3fe42;
               12'b000101010111: data1 <=  20'h01986;
               12'b000101011000: data1 <=  20'h028c9;
               12'b000101011001: data1 <=  20'h020c9;
               12'b000101011010: data1 <=  20'h4ed26;
               12'b000101011011: data1 <=  20'h265a6;
               12'b000101011100: data1 <=  20'h4ed26;
               12'b000101011101: data1 <=  20'h1fccf;
               12'b000101011110: data1 <=  20'h34126;
               12'b000101011111: data1 <=  20'h2786e;
               12'b000101100000: data1 <=  20'h4ed26;
               12'b000101100001: data1 <=  20'h4c144;
               12'b000101100010: data1 <=  20'h09893;
               12'b000101100011: data1 <=  20'h08093;
               12'b000101100100: data1 <=  20'h3ccc9;
               12'b000101100101: data1 <=  20'h83a43;
               12'b000101100110: data1 <=  20'h54d49;
               12'b000101100111: data1 <=  20'h51ac4;
               12'b000101101000: data1 <=  20'h26a06;
               12'b000101101001: data1 <=  20'h00656;
               12'b000101101010: data1 <=  20'h2e50e;
               12'b000101101011: data1 <=  20'h190d4;
               12'b000101101100: data1 <=  20'h03cc9;
               12'b000101101101: data1 <=  20'h00cc9;
               12'b000101101110: data1 <=  20'h4eccc;
               12'b000101101111: data1 <=  20'h4bccc;
               12'b000101110000: data1 <=  20'h4ed26;
               12'b000101110001: data1 <=  20'h4b126;
               12'b000101110010: data1 <=  20'h58a63;
               12'b000101110011: data1 <=  20'h51e63;
               12'b000101110100: data1 <=  20'h61546;
               12'b000101110101: data1 <=  20'h0194c;
               12'b000101110110: data1 <=  20'h0a8cc;
               12'b000101110111: data1 <=  20'h068cc;
               12'b000101111000: data1 <=  20'h5b8c9;
               12'b000101111001: data1 <=  20'h1492c;
               12'b000101111010: data1 <=  20'h0948c;
               12'b000101111011: data1 <=  20'h011c8;
               12'b000101111100: data1 <=  20'h280c9;
               12'b000101111101: data1 <=  20'h3f243;
               12'b000101111110: data1 <=  20'h61926;
               12'b000101111111: data1 <=  20'h066b7;
               12'b000110000000: data1 <=  20'h39e24;
               12'b000110000001: data1 <=  20'h00572;
               12'b000110000010: data1 <=  20'h5f5a6;
               12'b000110000011: data1 <=  20'h5dd26;
               12'b000110000100: data1 <=  20'h2dde4;
               12'b000110000101: data1 <=  20'h4d4c9;
               12'b000110000110: data1 <=  20'h33a43;
               12'b000110000111: data1 <=  20'h57b04;
               12'b000110001000: data1 <=  20'h4286c;
               12'b000110001001: data1 <=  20'h12f03;
               12'b000110001010: data1 <=  20'h6dd46;
               12'b000110001011: data1 <=  20'h51a43;
               12'b000110001100: data1 <=  20'h01649;
               12'b000110001101: data1 <=  20'h13e09;
               12'b000110001110: data1 <=  20'h2346c;
               12'b000110001111: data1 <=  20'h2be44;
               12'b000110010000: data1 <=  20'h280c9;
               12'b000110010001: data1 <=  20'h344ca;
               12'b000110010010: data1 <=  20'h600c9;
               12'b000110010011: data1 <=  20'h07255;
               12'b000110010100: data1 <=  20'h33987;
               12'b000110010101: data1 <=  20'h214c9;
               12'b000110010110: data1 <=  20'h0cb04;
               12'b000110010111: data1 <=  20'h2f4ac;
               12'b000110011000: data1 <=  20'h2d0ac;
               12'b000110011001: data1 <=  20'h27cc9;
               12'b000110011010: data1 <=  20'h064d1;
               12'b000110011011: data1 <=  20'h07269;
               12'b000110011100: data1 <=  20'h71586;
               12'b000110011101: data1 <=  20'h1e093;
               12'b000110011110: data1 <=  20'h64147;
               12'b000110011111: data1 <=  20'h2dd4c;
               12'b000110100000: data1 <=  20'h2d54c;
               12'b000110100001: data1 <=  20'h0ed26;
               12'b000110100010: data1 <=  20'h7d6a4;
               12'b000110100011: data1 <=  20'h4d526;
               12'b000110100100: data1 <=  20'h0e526;
               12'b000110100101: data1 <=  20'h0348e;
               12'b000110100110: data1 <=  20'h01c8e;
               12'b000110100111: data1 <=  20'h61526;
               12'b000110101000: data1 <=  20'h32a45;
               12'b000110101001: data1 <=  20'h174cb;
               12'b000110101010: data1 <=  20'h20d6e;
               12'b000110101011: data1 <=  20'h1d8c9;
               12'b000110101100: data1 <=  20'h27526;
               12'b000110101101: data1 <=  20'h1d8c9;
               12'b000110101110: data1 <=  20'h190c9;
               12'b000110101111: data1 <=  20'h1b524;
               12'b000110110000: data1 <=  20'h89a62;
               12'b000110110001: data1 <=  20'h5bcc9;
               12'b000110110010: data1 <=  20'h57cc9;
               12'b000110110011: data1 <=  20'h48489;
               12'b000110110100: data1 <=  20'h46489;
               12'b000110110101: data1 <=  20'h39247;
               12'b000110110110: data1 <=  20'h4d4ca;
               12'b000110110111: data1 <=  20'h030c9;
               12'b000110111000: data1 <=  20'h018c9;
               12'b000110111001: data1 <=  20'h6be43;
               12'b000110111010: data1 <=  20'h6aa43;
               12'b000110111011: data1 <=  20'h2816c;
               12'b000110111100: data1 <=  20'h26dc6;
               12'b000110111101: data1 <=  20'h1a5e4;
               12'b000110111110: data1 <=  20'h002c2;
               12'b000110111111: data1 <=  20'h00318;
               12'b000111000000: data1 <=  20'h5e244;
               12'b000111000001: data1 <=  20'h33989;
               12'b000111000010: data1 <=  20'h4c0ec;
               12'b000111000011: data1 <=  20'h0cec6;
               12'b000111000100: data1 <=  20'h7e5c3;
               12'b000111000101: data1 <=  20'h00310;
               12'b000111000110: data1 <=  20'h52244;
               12'b000111000111: data1 <=  20'h3f2c2;
               12'b000111001000: data1 <=  20'h14568;
               12'b000111001001: data1 <=  20'h22cc6;
               12'b000111001010: data1 <=  20'h2bf06;
               12'b000111001011: data1 <=  20'h0394a;
               12'b000111001100: data1 <=  20'h0014a;
               12'b000111001101: data1 <=  20'h06704;
               12'b000111001110: data1 <=  20'h6a643;
               12'b000111001111: data1 <=  20'h5f206;
               12'b000111010000: data1 <=  20'h5ea06;
               12'b000111010001: data1 <=  20'h65a43;
               12'b000111010010: data1 <=  20'h516aa;
               12'b000111010011: data1 <=  20'h034d8;
               12'b000111010100: data1 <=  20'h1accb;
               12'b000111010101: data1 <=  20'h21926;
               12'b000111010110: data1 <=  20'h19454;
               12'b000111010111: data1 <=  20'h034d8;
               12'b000111011000: data1 <=  20'h014d8;
               12'b000111011001: data1 <=  20'h2fcce;
               12'b000111011010: data1 <=  20'h2cc8c;
               12'b000111011011: data1 <=  20'h1f70e;
               12'b000111011100: data1 <=  20'h52946;
               12'b000111011101: data1 <=  20'h030c9;
               12'b000111011110: data1 <=  20'h2c4ce;
               12'b000111011111: data1 <=  20'h1052f;
               12'b000111100000: data1 <=  20'h0c8c9;
               12'b000111100001: data1 <=  20'h0f94e;
               12'b000111100010: data1 <=  20'h28452;
               12'b000111100011: data1 <=  20'h219e6;
               12'b000111100100: data1 <=  20'h278ca;
               12'b000111100101: data1 <=  20'h030c9;
               12'b000111100110: data1 <=  20'h13927;
               12'b000111100111: data1 <=  20'h2d5c3;
               12'b000111101000: data1 <=  20'h2d906;
               12'b000111101001: data1 <=  20'h2ecec;
               12'b000111101010: data1 <=  20'h28092;
               12'b000111101011: data1 <=  20'h5b8c9;
               12'b000111101100: data1 <=  20'h010cd;
               12'b000111101101: data1 <=  20'h0d2a3;
               12'b000111101110: data1 <=  20'h1a4ac;
               12'b000111101111: data1 <=  20'h1548a;
               12'b000111110000: data1 <=  20'h1b0a8;
               12'b000111110001: data1 <=  20'h01969;
               12'b000111110010: data1 <=  20'h27185;
               12'b000111110011: data1 <=  20'h00305;
               12'b000111110100: data1 <=  20'h3eee6;
               12'b000111110101: data1 <=  20'h84243;
               12'b000111110110: data1 <=  20'h266a6;
               12'b000111110111: data1 <=  20'h1f4cc;
               12'b000111111000: data1 <=  20'h0f08f;
               12'b000111111001: data1 <=  20'h2dd0a;
               12'b000111111010: data1 <=  20'h2d1ec;
               12'b000111111011: data1 <=  20'h6a546;
               12'b000111111100: data1 <=  20'h74126;
               12'b000111111101: data1 <=  20'h27cd0;
               12'b000111111110: data1 <=  20'h74126;
               12'b000111111111: data1 <=  20'h70d26;
               12'b001000000000: data1 <=  20'h3c126;
               12'b001000000001: data1 <=  20'h38526;
               12'b001000000010: data1 <=  20'h170c9;
               12'b001000000011: data1 <=  20'h6ae43;
               12'b001000000100: data1 <=  20'h5eaa6;
               12'b001000000101: data1 <=  20'h6c8c6;
               12'b001000000110: data1 <=  20'h174c9;
               12'b001000000111: data1 <=  20'h12cc9;
               12'b001000001000: data1 <=  20'h0120a;
               12'b001000001001: data1 <=  20'h00950;
               12'b001000001010: data1 <=  20'h03945;
               12'b001000001011: data1 <=  20'h00145;
               12'b001000001100: data1 <=  20'h174ca;
               12'b001000001101: data1 <=  20'h46186;
               12'b001000001110: data1 <=  20'h05472;
               12'b001000001111: data1 <=  20'h018c9;
               12'b001000010000: data1 <=  20'h34127;
               12'b001000010001: data1 <=  20'h4cd0a;
               12'b001000010010: data1 <=  20'h05472;
               12'b001000010011: data1 <=  20'h28089;
               12'b001000010100: data1 <=  20'h03d26;
               12'b001000010101: data1 <=  20'h0cb03;
               12'b001000010110: data1 <=  20'h2e8c9;
               12'b001000010111: data1 <=  20'h274ca;
               12'b001000011000: data1 <=  20'h094cc;
               12'b001000011001: data1 <=  20'h1a98c;
               12'b001000011010: data1 <=  20'h16455;
               12'b001000011011: data1 <=  20'h07d88;
               12'b001000011100: data1 <=  20'h00e48;
               12'b001000011101: data1 <=  20'h00e43;
               12'b001000011110: data1 <=  20'h51704;
               12'b001000011111: data1 <=  20'h21c89;
               12'b001000100000: data1 <=  20'h090c9;
               12'b001000100001: data1 <=  20'h0e0d6;
               12'b001000100010: data1 <=  20'h4290e;
               12'b001000100011: data1 <=  20'h19e0f;
               12'b001000100100: data1 <=  20'h4290e;
               12'b001000100101: data1 <=  20'h3e90e;
               12'b001000100110: data1 <=  20'h5a166;
               12'b001000100111: data1 <=  20'h2bf09;
               12'b001000101000: data1 <=  20'h09890;
               12'b001000101001: data1 <=  20'h08090;
               12'b001000101010: data1 <=  20'h20a08;
               12'b001000101011: data1 <=  20'h384c9;
               12'b001000101100: data1 <=  20'h65a43;
               12'b001000101101: data1 <=  20'h4bcc9;
               12'b001000101110: data1 <=  20'h59926;
               12'b001000101111: data1 <=  20'h51d0a;
               12'b001000110000: data1 <=  20'h23072;
               12'b001000110001: data1 <=  20'h20243;
               12'b001000110010: data1 <=  20'h238cb;
               12'b001000110011: data1 <=  20'h1f8cb;
               12'b001000110100: data1 <=  20'h0b089;
               12'b001000110101: data1 <=  20'h06889;
               12'b001000110110: data1 <=  20'h5ee49;
               12'b001000110111: data1 <=  20'h39d84;
               12'b001000111000: data1 <=  20'h10526;
               12'b001000111001: data1 <=  20'h0c926;
               12'b001000111010: data1 <=  20'h03cd1;
               12'b001000111011: data1 <=  20'h00cd1;
               12'b001000111100: data1 <=  20'h6c524;
               12'b001000111101: data1 <=  20'h20c72;
               12'b001000111110: data1 <=  20'h0ddcc;
               12'b001000111111: data1 <=  20'h0f06c;
               12'b001001000000: data1 <=  20'h2e5cf;
               12'b001001000001: data1 <=  20'h2bdcf;
               12'b001001000010: data1 <=  20'h03d26;
               12'b001001000011: data1 <=  20'h00126;
               12'b001001000100: data1 <=  20'h288ce;
               12'b001001000101: data1 <=  20'h2e0c9;
               12'b001001000110: data1 <=  20'h288cf;
               12'b001001000111: data1 <=  20'h270cf;
               12'b001001001000: data1 <=  20'h16909;
               12'b001001001001: data1 <=  20'h00135;
               12'b001001001010: data1 <=  20'h3b10c;
               12'b001001001011: data1 <=  20'h2d54c;
               12'b001001001100: data1 <=  20'h28092;
               12'b001001001101: data1 <=  20'h000c9;
               12'b001001001110: data1 <=  20'h58643;
               12'b001001001111: data1 <=  20'h5850a;
               12'b001001010000: data1 <=  20'h4b304;
               12'b001001010001: data1 <=  20'h0c874;
               12'b001001010010: data1 <=  20'h67148;
               12'b001001010011: data1 <=  20'h64948;
               12'b001001010100: data1 <=  20'h01d49;
               12'b001001010101: data1 <=  20'h00303;
               12'b001001010110: data1 <=  20'h32de4;
               12'b001001010111: data1 <=  20'h20d86;
               12'b001001011000: data1 <=  20'h529c6;
               12'b001001011001: data1 <=  20'h5a48a;
               12'b001001011010: data1 <=  20'h258c7;
               12'b001001011011: data1 <=  20'h048c6;
               12'b001001011100: data1 <=  20'h07243;
               12'b001001011101: data1 <=  20'h27dd2;
               12'b001001011110: data1 <=  20'h000c6;
               12'b001001011111: data1 <=  20'h480c6;
               12'b001001100000: data1 <=  20'h7d303;
               12'b001001100001: data1 <=  20'h480c7;
               12'b001001100010: data1 <=  20'h4c146;
               12'b001001100011: data1 <=  20'h480c6;
               12'b001001100100: data1 <=  20'h460c7;
               12'b001001100101: data1 <=  20'h1ad6c;
               12'b001001100110: data1 <=  20'h5f544;
               12'b001001100111: data1 <=  20'h038c9;
               12'b001001101000: data1 <=  20'h010c9;
               12'b001001101001: data1 <=  20'h0f48f;
               12'b001001101010: data1 <=  20'h00283;
               12'b001001101011: data1 <=  20'h73d46;
               12'b001001101100: data1 <=  20'h2c4cb;
               12'b001001101101: data1 <=  20'h5a149;
               12'b001001101110: data1 <=  20'h0e889;
               12'b001001101111: data1 <=  20'h16544;
               12'b001001110000: data1 <=  20'h27186;
               12'b001001110001: data1 <=  20'h3410a;
               12'b001001110010: data1 <=  20'h1ac90;
               12'b001001110011: data1 <=  20'h34124;
               12'b001001110100: data1 <=  20'h0ddc9;
               12'b001001110101: data1 <=  20'h64e68;
               12'b001001110110: data1 <=  20'h00148;
               12'b001001110111: data1 <=  20'h0de12;
               12'b001001111000: data1 <=  20'h44f0b;
               12'b001001111001: data1 <=  20'h13a45;
               12'b001001111010: data1 <=  20'h64643;
               12'b001001111011: data1 <=  20'h6ba43;
               12'b001001111100: data1 <=  20'h51926;
               12'b001001111101: data1 <=  20'h38aea;
               12'b001001111110: data1 <=  20'h2ca43;
               12'b001001111111: data1 <=  20'h33983;
               12'b001010000000: data1 <=  20'h0e076;
               12'b001010000001: data1 <=  20'h6dd46;
               12'b001010000010: data1 <=  20'h70d46;
               12'b001010000011: data1 <=  20'h158cc;
               12'b001010000100: data1 <=  20'h28089;
               12'b001010000101: data1 <=  20'h02cc9;
               12'b001010000110: data1 <=  20'h01cc9;
               12'b001010000111: data1 <=  20'h41926;
               12'b001010001000: data1 <=  20'h454c9;
               12'b001010001001: data1 <=  20'h22c73;
               12'b001010001010: data1 <=  20'h27126;
               12'b001010001011: data1 <=  20'h22c73;
               12'b001010001100: data1 <=  20'h12cc9;
               12'b001010001101: data1 <=  20'h84a43;
               12'b001010001110: data1 <=  20'h3ee44;
               12'b001010001111: data1 <=  20'h1c50a;
               12'b001010010000: data1 <=  20'h33d26;
               12'b001010010001: data1 <=  20'h3b528;
               12'b001010010010: data1 <=  20'h258ac;
               12'b001010010011: data1 <=  20'h275c6;
               12'b001010010100: data1 <=  20'h21073;
               12'b001010010101: data1 <=  20'h1b1f4;
               12'b001010010110: data1 <=  20'h195f4;
               12'b001010010111: data1 <=  20'h41cc6;
               12'b001010011000: data1 <=  20'h3fcc6;
               12'b001010011001: data1 <=  20'h100ce;
               12'b001010011010: data1 <=  20'h0d8ce;
               12'b001010011011: data1 <=  20'h1c0c7;
               12'b001010011100: data1 <=  20'h1b4c9;
               12'b001010011101: data1 <=  20'h1bd0a;
               12'b001010011110: data1 <=  20'h1a50a;
               12'b001010011111: data1 <=  20'h72946;
               12'b001010100000: data1 <=  20'h70ea6;
               12'b001010100001: data1 <=  20'h0ed86;
               12'b001010100010: data1 <=  20'h0d586;
               12'b001010100011: data1 <=  20'h22586;
               12'b001010100100: data1 <=  20'h340c9;
               12'b001010100101: data1 <=  20'h2c686;
               12'b001010100110: data1 <=  20'h1f586;
               12'b001010100111: data1 <=  20'h5b10a;
               12'b001010101000: data1 <=  20'h5810a;
               12'b001010101001: data1 <=  20'h4568d;
               12'b001010101010: data1 <=  20'h39d85;
               12'b001010101011: data1 <=  20'h26e06;
               12'b001010101100: data1 <=  20'h77124;
               12'b001010101101: data1 <=  20'h21185;
               12'b001010101110: data1 <=  20'h201cc;
               12'b001010101111: data1 <=  20'h1b526;
               12'b001010110000: data1 <=  20'h26263;
               12'b001010110001: data1 <=  20'h430c9;
               12'b001010110010: data1 <=  20'h2ca42;
               12'b001010110011: data1 <=  20'h11892;
               12'b001010110100: data1 <=  20'h71283;
               12'b001010110101: data1 <=  20'h38ac3;
               12'b001010110110: data1 <=  20'h0c892;
               12'b001010110111: data1 <=  20'h04c97;
               12'b001010111000: data1 <=  20'h12cd3;
               12'b001010111001: data1 <=  20'h110c9;
               12'b001010111010: data1 <=  20'h1f546;
               12'b001010111011: data1 <=  20'h01d8c;
               12'b001010111100: data1 <=  20'h12f06;
               12'b001010111101: data1 <=  20'h5a08a;
               12'b001010111110: data1 <=  20'h3a48f;
               12'b001010111111: data1 <=  20'h45e26;
               12'b001011000000: data1 <=  20'h1fe48;
               12'b001011000001: data1 <=  20'h275c6;
               12'b001011000010: data1 <=  20'h265c6;
               12'b001011000011: data1 <=  20'h23472;
               12'b001011000100: data1 <=  20'h20872;
               12'b001011000101: data1 <=  20'h411c4;
               12'b001011000110: data1 <=  20'h3f924;
               12'b001011000111: data1 <=  20'h00a49;
               12'b001011001000: data1 <=  20'h14588;
               12'b001011001001: data1 <=  20'h06905;
               12'b001011001010: data1 <=  20'h2ece8;
               12'b001011001011: data1 <=  20'h4b2c4;
               12'b001011001100: data1 <=  20'h2948f;
               12'b001011001101: data1 <=  20'h2d0e8;
               12'b001011001110: data1 <=  20'h72924;
               12'b001011001111: data1 <=  20'h0cec4;
               12'b001011010000: data1 <=  20'h170d1;
               12'b001011010001: data1 <=  20'h0e912;
               12'b001011010010: data1 <=  20'h044cc;
               12'b001011010011: data1 <=  20'h01cc9;
               12'b001011010100: data1 <=  20'h2312c;
               12'b001011010101: data1 <=  20'h8a242;
               12'b001011010110: data1 <=  20'h41186;
               12'b001011010111: data1 <=  20'h0648b;
               12'b001011011000: data1 <=  20'h0508a;
               12'b001011011001: data1 <=  20'h130d1;
               12'b001011011010: data1 <=  20'h61926;
               12'b001011011011: data1 <=  20'h51509;
               12'b001011011100: data1 <=  20'h360cc;
               12'b001011011101: data1 <=  20'h328cc;
               12'b001011011110: data1 <=  20'h0f08f;
               12'b001011011111: data1 <=  20'h1fa63;
               12'b001011100000: data1 <=  20'h34d27;
               12'b001011100001: data1 <=  20'h32d89;
               12'b001011100010: data1 <=  20'h26643;
               12'b001011100011: data1 <=  20'h0288c;
               12'b001011100100: data1 <=  20'h3924e;
               12'b001011100101: data1 <=  20'h00089;
               12'b001011100110: data1 <=  20'h22492;
               12'b001011100111: data1 <=  20'h21492;
               12'b001011101000: data1 <=  20'h21cca;
               12'b001011101001: data1 <=  20'h1b48b;
               12'b001011101010: data1 <=  20'h65243;
               12'b001011101011: data1 <=  20'h64283;
               12'b001011101100: data1 <=  20'h3a8cc;
               12'b001011101101: data1 <=  20'h53508;
               12'b001011101110: data1 <=  20'h41c6c;
               12'b001011101111: data1 <=  20'h399ce;
               12'b001011110000: data1 <=  20'h0030a;
               12'b001011110001: data1 <=  20'h45242;
               12'b001011110010: data1 <=  20'h240ac;
               12'b001011110011: data1 <=  20'h1f4ac;
               12'b001011110100: data1 <=  20'h29912;
               12'b001011110101: data1 <=  20'h25912;
               12'b001011110110: data1 <=  20'h2258c;
               12'b001011110111: data1 <=  20'h274c9;
               12'b001011111000: data1 <=  20'h538cb;
               12'b001011111001: data1 <=  20'h1f58c;
               12'b001011111010: data1 <=  20'h0cee3;
               12'b001011111011: data1 <=  20'h5e263;
               12'b001011111100: data1 <=  20'h6d964;
               12'b001011111101: data1 <=  20'h51505;
               12'b001011111110: data1 <=  20'h41944;
               12'b001011111111: data1 <=  20'h26929;
               12'b001100000000: data1 <=  20'h5b526;
               12'b001100000001: data1 <=  20'h4b526;
               12'b001100000010: data1 <=  20'h3f688;
               12'b001100000011: data1 <=  20'h00932;
               12'b001100000100: data1 <=  20'h4812a;
               12'b001100000101: data1 <=  20'h0cd05;
               12'b001100000110: data1 <=  20'h19ea6;
               12'b001100000111: data1 <=  20'h01d4e;
               12'b001100001000: data1 <=  20'h6d584;
               12'b001100001001: data1 <=  20'h25ae4;
               12'b001100001010: data1 <=  20'h41d0a;
               12'b001100001011: data1 <=  20'h64243;
               12'b001100001100: data1 <=  20'h67d24;
               12'b001100001101: data1 <=  20'h64124;
               12'b001100001110: data1 <=  20'h480c6;
               12'b001100001111: data1 <=  20'h460c6;
               12'b001100010000: data1 <=  20'h12f06;
               12'b001100010001: data1 <=  20'h19a43;
               12'b001100010010: data1 <=  20'h00304;
               12'b001100010011: data1 <=  20'h64643;
               12'b001100010100: data1 <=  20'h61926;
               12'b001100010101: data1 <=  20'h5dd26;
               12'b001100010110: data1 <=  20'h6be43;
               12'b001100010111: data1 <=  20'h340ca;
               12'b001100011000: data1 <=  20'h280c9;
               12'b001100011001: data1 <=  20'h340a8;
               12'b001100011010: data1 <=  20'h350c8;
               12'b001100011011: data1 <=  20'h20ccb;
               12'b001100011100: data1 <=  20'h28d09;
               12'b001100011101: data1 <=  20'h2c2a6;
               12'b001100011110: data1 <=  20'h2306c;
               12'b001100011111: data1 <=  20'h39d6c;
               12'b001100100000: data1 <=  20'h35548;
               12'b001100100001: data1 <=  20'h33583;
               12'b001100100010: data1 <=  20'h46644;
               12'b001100100011: data1 <=  20'h002d6;
               12'b001100100100: data1 <=  20'h0f4c8;
               12'b001100100101: data1 <=  20'h024c9;
               12'b001100100110: data1 <=  20'h028c9;
               12'b001100100111: data1 <=  20'h14cce;
               12'b001100101000: data1 <=  20'h3f648;
               12'b001100101001: data1 <=  20'h0286e;
               12'b001100101010: data1 <=  20'h13e14;
               12'b001100101011: data1 <=  20'h1b4ca;
               12'b001100101100: data1 <=  20'h01604;
               12'b001100101101: data1 <=  20'h1fe44;
               12'b001100101110: data1 <=  20'h034c9;
               12'b001100101111: data1 <=  20'h1b105;
               12'b001100110000: data1 <=  20'h41944;
               12'b001100110001: data1 <=  20'h3f144;
               12'b001100110010: data1 <=  20'h46985;
               12'b001100110011: data1 <=  20'h3f50a;
               12'b001100110100: data1 <=  20'h4dd28;
               12'b001100110101: data1 <=  20'h83703;
               12'b001100110110: data1 <=  20'h7de44;
               12'b001100110111: data1 <=  20'h5e126;
               12'b001100111000: data1 <=  20'h6d144;
               12'b001100111001: data1 <=  20'h4d48c;
               12'b001100111010: data1 <=  20'h27d26;
               12'b001100111011: data1 <=  20'h518c9;
               12'b001100111100: data1 <=  20'h65984;
               12'b001100111101: data1 <=  20'h1fa83;
               12'b001100111110: data1 <=  20'h08529;
               12'b001100111111: data1 <=  20'h77524;
               12'b001101000000: data1 <=  20'h09092;
               12'b001101000001: data1 <=  20'h0e50c;
               12'b001101000010: data1 <=  20'h41528;
               12'b001101000011: data1 <=  20'h46185;
               12'b001101000100: data1 <=  20'h3b126;
               12'b001101000101: data1 <=  20'h3fcc9;
               12'b001101000110: data1 <=  20'h2ccac;
               12'b001101000111: data1 <=  20'h00aa6;
               12'b001101001000: data1 <=  20'h27546;
               12'b001101001001: data1 <=  20'h024cf;
               12'b001101001010: data1 <=  20'h0d242;
               12'b001101001011: data1 <=  20'h6c506;
               12'b001101001100: data1 <=  20'h00e42;
               12'b001101001101: data1 <=  20'h02126;
               12'b001101001110: data1 <=  20'h6a643;
               12'b001101001111: data1 <=  20'h2d585;
               12'b001101010000: data1 <=  20'h12cc9;
               12'b001101010001: data1 <=  20'h11889;
               12'b001101010010: data1 <=  20'h0c889;
               12'b001101010011: data1 <=  20'h06704;
               12'b001101010100: data1 <=  20'h64126;
               12'b001101010101: data1 <=  20'h54d26;
               12'b001101010110: data1 <=  20'h5de63;
               12'b001101010111: data1 <=  20'h1facc;
               12'b001101011000: data1 <=  20'h528c6;
               12'b001101011001: data1 <=  20'h0da83;
               12'b001101011010: data1 <=  20'h598ca;
               12'b001101011011: data1 <=  20'h4ca06;
               12'b001101011100: data1 <=  20'h51d09;
               12'b001101011101: data1 <=  20'h34cce;
               12'b001101011110: data1 <=  20'h4ba06;
               12'b001101011111: data1 <=  20'h65608;
               12'b001101100000: data1 <=  20'h0888c;
               12'b001101100001: data1 <=  20'h0e90a;
               12'b001101100010: data1 <=  20'h27186;
               12'b001101100011: data1 <=  20'h2e4c9;
               12'b001101100100: data1 <=  20'h0010c;
               12'b001101100101: data1 <=  20'h368c9;
               12'b001101100110: data1 <=  20'h4b8c6;
               12'b001101100111: data1 <=  20'h842a3;
               12'b001101101000: data1 <=  20'h00a06;
               12'b001101101001: data1 <=  20'h28ce6;
               12'b001101101010: data1 <=  20'h1a88e;
               12'b001101101011: data1 <=  20'h2e0c9;
               12'b001101101100: data1 <=  20'h33cce;
               12'b001101101101: data1 <=  20'h36890;
               12'b001101101110: data1 <=  20'h59cca;
               12'b001101101111: data1 <=  20'h46585;
               12'b001101110000: data1 <=  20'h4b2e3;
               12'b001101110001: data1 <=  20'h034cc;
               12'b001101110010: data1 <=  20'h3e985;
               12'b001101110011: data1 <=  20'h0fd44;
               12'b001101110100: data1 <=  20'h014cc;
               12'b001101110101: data1 <=  20'h28526;
               12'b001101110110: data1 <=  20'h26926;
               12'b001101110111: data1 <=  20'h4664d;
               12'b001101111000: data1 <=  20'h44e4d;
               12'b001101111001: data1 <=  20'h67186;
               12'b001101111010: data1 <=  20'h25aa3;
               12'b001101111011: data1 <=  20'h67186;
               12'b001101111100: data1 <=  20'h2d0ce;
               12'b001101111101: data1 <=  20'h3fe62;
               12'b001101111110: data1 <=  20'h1a5c4;
               12'b001101111111: data1 <=  20'h71644;
               12'b001110000000: data1 <=  20'h01c89;
               12'b001110000001: data1 <=  20'h16164;
               12'b001110000010: data1 <=  20'h00926;
               12'b001110000011: data1 <=  20'h0b097;
               12'b001110000100: data1 <=  20'h06897;
               12'b001110000101: data1 <=  20'h65643;
               12'b001110000110: data1 <=  20'h12d64;
               12'b001110000111: data1 <=  20'h64a83;
               12'b001110001000: data1 <=  20'h141a4;
               12'b001110001001: data1 <=  20'h38acf;
               12'b001110001010: data1 <=  20'h19dc3;
               12'b001110001011: data1 <=  20'h2dd44;
               12'b001110001100: data1 <=  20'h2d544;
               12'b001110001101: data1 <=  20'h1b8c9;
               12'b001110001110: data1 <=  20'h4b526;
               12'b001110001111: data1 <=  20'h14d0a;
               12'b001110010000: data1 <=  20'h26606;
               12'b001110010001: data1 <=  20'h26dc6;
               12'b001110010010: data1 <=  20'h13d26;
               12'b001110010011: data1 <=  20'h14642;
               12'b001110010100: data1 <=  20'h27526;
               12'b001110010101: data1 <=  20'h06703;
               12'b001110010110: data1 <=  20'h6a546;
               12'b001110010111: data1 <=  20'h71643;
               12'b001110011000: data1 <=  20'h1fcd0;
               12'b001110011001: data1 <=  20'h27566;
               12'b001110011010: data1 <=  20'h0dd96;
               12'b001110011011: data1 <=  20'h2e48a;
               12'b001110011100: data1 <=  20'h02492;
               12'b001110011101: data1 <=  20'h368c9;
               12'b001110011110: data1 <=  20'h2cdea;
               12'b001110011111: data1 <=  20'h21cc9;
               12'b001110100000: data1 <=  20'h3a8ca;
               12'b001110100001: data1 <=  20'h5a4ca;
               12'b001110100010: data1 <=  20'h594ca;
               12'b001110100011: data1 <=  20'h33209;
               12'b001110100100: data1 <=  20'h45683;
               12'b001110100101: data1 <=  20'h0348d;
               12'b001110100110: data1 <=  20'h01c8d;
               12'b001110100111: data1 <=  20'h07247;
               12'b001110101000: data1 <=  20'h450c9;
               12'b001110101001: data1 <=  20'h72926;
               12'b001110101010: data1 <=  20'h391e6;
               12'b001110101011: data1 <=  20'h3fe62;
               12'b001110101100: data1 <=  20'h278f0;
               12'b001110101101: data1 <=  20'h59d26;
               12'b001110101110: data1 <=  20'h2bd0c;
               12'b001110101111: data1 <=  20'h1aa43;
               12'b001110110000: data1 <=  20'h64186;
               12'b001110110001: data1 <=  20'h54924;
               12'b001110110010: data1 <=  20'h335ce;
               12'b001110110011: data1 <=  20'h646c6;
               12'b001110110100: data1 <=  20'h024c9;
               12'b001110110101: data1 <=  20'h2194a;
               12'b001110110110: data1 <=  20'h2094a;
               12'b001110110111: data1 <=  20'h26a06;
               12'b001110111000: data1 <=  20'h2bcc9;
               12'b001110111001: data1 <=  20'h4290e;
               12'b001110111010: data1 <=  20'h4d4cc;
               12'b001110111011: data1 <=  20'h4090c;
               12'b001110111100: data1 <=  20'h02089;
               12'b001110111101: data1 <=  20'h1b910;
               12'b001110111110: data1 <=  20'h40546;
               12'b001110111111: data1 <=  20'h26dce;
               12'b001111000000: data1 <=  20'h45682;
               12'b001111000001: data1 <=  20'h36890;
               12'b001111000010: data1 <=  20'h4518a;
               12'b001111000011: data1 <=  20'h39d84;
               12'b001111000100: data1 <=  20'h4d4c7;
               12'b001111000101: data1 <=  20'h1b910;
               12'b001111000110: data1 <=  20'h1a910;
               12'b001111000111: data1 <=  20'h3a526;
               12'b001111001000: data1 <=  20'h1fa0c;
               12'b001111001001: data1 <=  20'h3a8c8;
               12'b001111001010: data1 <=  20'h01872;
               12'b001111001011: data1 <=  20'h3c8ae;
               12'b001111001100: data1 <=  20'h38cae;
               12'b001111001101: data1 <=  20'h1ad46;
               12'b001111001110: data1 <=  20'h132f2;
               12'b001111001111: data1 <=  20'h06aa3;
               12'b001111010000: data1 <=  20'h27cc9;
               12'b001111010001: data1 <=  20'h71586;
               12'b001111010010: data1 <=  20'h36110;
               12'b001111010011: data1 <=  20'h76f04;
               12'b001111010100: data1 <=  20'h36110;
               12'b001111010101: data1 <=  20'h32110;
               12'b001111010110: data1 <=  20'h4d10a;
               12'b001111010111: data1 <=  20'h2d0a8;
               12'b001111011000: data1 <=  20'h07662;
               12'b001111011001: data1 <=  20'h4b309;
               12'b001111011010: data1 <=  20'h019a8;
               12'b001111011011: data1 <=  20'h00303;
               12'b001111011100: data1 <=  20'h17c8b;
               12'b001111011101: data1 <=  20'h278c9;
               12'b001111011110: data1 <=  20'h46588;
               12'b001111011111: data1 <=  20'h32186;
               12'b001111100000: data1 <=  20'h6be43;
               12'b001111100001: data1 <=  20'h57926;
               12'b001111100010: data1 <=  20'h17c89;
               12'b001111100011: data1 <=  20'h12c89;
               12'b001111100100: data1 <=  20'h03d33;
               12'b001111100101: data1 <=  20'h00133;
               12'b001111100110: data1 <=  20'h480c8;
               12'b001111100111: data1 <=  20'h460c8;
               12'b001111101000: data1 <=  20'h46263;
               12'b001111101001: data1 <=  20'h7de44;
               12'b001111101010: data1 <=  20'h27206;
               12'b001111101011: data1 <=  20'h01926;
               12'b001111101100: data1 <=  20'h1548e;
               12'b001111101101: data1 <=  20'h1f9ec;
               12'b001111101110: data1 <=  20'h4dd05;
               12'b001111101111: data1 <=  20'h014c9;
               12'b001111110000: data1 <=  20'h030c9;
               12'b001111110001: data1 <=  20'h20988;
               12'b001111110010: data1 <=  20'h4e566;
               12'b001111110011: data1 <=  20'h516a3;
               12'b001111110100: data1 <=  20'h0850c;
               12'b001111110101: data1 <=  20'h004cc;
               12'b001111110110: data1 <=  20'h0d2a2;
               12'b001111110111: data1 <=  20'h0d263;
               12'b001111111000: data1 <=  20'h42cce;
               12'b001111111001: data1 <=  20'h3ecce;
               12'b001111111010: data1 <=  20'h275ce;
               12'b001111111011: data1 <=  20'h4b126;
               12'b001111111100: data1 <=  20'h5b509;
               12'b001111111101: data1 <=  20'h06ac4;
               12'b001111111110: data1 <=  20'h47126;
               12'b001111111111: data1 <=  20'h5de43;
               12'b010000000000: data1 <=  20'h5b8e9;
               12'b010000000001: data1 <=  20'h13e04;
               12'b010000000010: data1 <=  20'h27585;
               12'b010000000011: data1 <=  20'h27c89;
               12'b010000000100: data1 <=  20'h0948a;
               12'b010000000101: data1 <=  20'h0848a;
               12'b010000000110: data1 <=  20'h618c9;
               12'b010000000111: data1 <=  20'h5e8c9;
               12'b010000001000: data1 <=  20'h0a073;
               12'b010000001001: data1 <=  20'h130c9;
               12'b010000001010: data1 <=  20'h03c73;
               12'b010000001011: data1 <=  20'h14584;
               12'b010000001100: data1 <=  20'h21c89;
               12'b010000001101: data1 <=  20'h01873;
               12'b010000001110: data1 <=  20'h0906c;
               12'b010000001111: data1 <=  20'h2d545;
               12'b010000010000: data1 <=  20'h15872;
               12'b010000010001: data1 <=  20'h150cc;
               12'b010000010010: data1 <=  20'h2ca63;
               12'b010000010011: data1 <=  20'h2c643;
               12'b010000010100: data1 <=  20'h52244;
               12'b010000010101: data1 <=  20'h200c9;
               12'b010000010110: data1 <=  20'h07684;
               12'b010000010111: data1 <=  20'h06684;
               12'b010000011000: data1 <=  20'h604c6;
               12'b010000011001: data1 <=  20'h0cb08;
               12'b010000011010: data1 <=  20'h20a43;
               12'b010000011011: data1 <=  20'h5fcc6;
               12'b010000011100: data1 <=  20'h4dd05;
               12'b010000011101: data1 <=  20'h4c505;
               12'b010000011110: data1 <=  20'h015c6;
               12'b010000011111: data1 <=  20'h0f08f;
               12'b010000100000: data1 <=  20'h2e4ac;
               12'b010000100001: data1 <=  20'h3a10e;
               12'b010000100010: data1 <=  20'h1fac6;
               12'b010000100011: data1 <=  20'h1f4c6;
               12'b010000100100: data1 <=  20'h6d524;
               12'b010000100101: data1 <=  20'h71263;
               12'b010000100110: data1 <=  20'h6d524;
               12'b010000100111: data1 <=  20'h6aa43;
               12'b010000101000: data1 <=  20'h6d524;
               12'b010000101001: data1 <=  20'h00303;
               12'b010000101010: data1 <=  20'h015c4;
               12'b010000101011: data1 <=  20'h59126;
               12'b010000101100: data1 <=  20'h54cc9;
               12'b010000101101: data1 <=  20'h7e5a4;
               12'b010000101110: data1 <=  20'h3a8cc;
               12'b010000101111: data1 <=  20'h3eea3;
               12'b010000110000: data1 <=  20'h34126;
               12'b010000110001: data1 <=  20'h3f527;
               12'b010000110010: data1 <=  20'h41948;
               12'b010000110011: data1 <=  20'h5df03;
               12'b010000110100: data1 <=  20'h21526;
               12'b010000110101: data1 <=  20'h524c9;
               12'b010000110110: data1 <=  20'h6d524;
               12'b010000110111: data1 <=  20'h4d4c6;
               12'b010000111000: data1 <=  20'h3a9ca;
               12'b010000111001: data1 <=  20'h389ca;
               12'b010000111010: data1 <=  20'h2dd31;
               12'b010000111011: data1 <=  20'h19cd4;
               12'b010000111100: data1 <=  20'h33d44;
               12'b010000111101: data1 <=  20'h2e489;
               12'b010000111110: data1 <=  20'h604c9;
               12'b010000111111: data1 <=  20'h32cd0;
               12'b010001000000: data1 <=  20'h6d524;
               12'b010001000001: data1 <=  20'h6b124;
               12'b010001000010: data1 <=  20'h08d26;
               12'b010001000011: data1 <=  20'h2d08a;
               12'b010001000100: data1 <=  20'h21186;
               12'b010001000101: data1 <=  20'h1a928;
               12'b010001000110: data1 <=  20'h67148;
               12'b010001000111: data1 <=  20'h64948;
               12'b010001001000: data1 <=  20'h00304;
               12'b010001001001: data1 <=  20'h25926;
               12'b010001001010: data1 <=  20'h19306;
               12'b010001001011: data1 <=  20'h01564;
               12'b010001001100: data1 <=  20'h06ac4;
               12'b010001001101: data1 <=  20'h27cd2;
               12'b010001001110: data1 <=  20'h38e84;
               12'b010001001111: data1 <=  20'h0ddce;
               12'b010001010000: data1 <=  20'h0da06;
               12'b010001010001: data1 <=  20'h13663;
               12'b010001010010: data1 <=  20'h08144;
               12'b010001010011: data1 <=  20'h3848f;
               12'b010001010100: data1 <=  20'h3f2a3;
               12'b010001010101: data1 <=  20'h00cc6;
               12'b010001010110: data1 <=  20'h1a9c9;
               12'b010001010111: data1 <=  20'h088c9;
               12'b010001011000: data1 <=  20'h35d29;
               12'b010001011001: data1 <=  20'h02095;
               12'b010001011010: data1 <=  20'h8a662;
               12'b010001011011: data1 <=  20'h5e683;
               12'b010001011100: data1 <=  20'h04c8d;
               12'b010001011101: data1 <=  20'h2c108;
               12'b010001011110: data1 <=  20'h5b0c9;
               12'b010001011111: data1 <=  20'h588c9;
               12'b010001100000: data1 <=  20'h22c8a;
               12'b010001100001: data1 <=  20'h20c8a;
               12'b010001100010: data1 <=  20'h22cc6;
               12'b010001100011: data1 <=  20'h204c6;
               12'b010001100100: data1 <=  20'h0cb15;
               12'b010001100101: data1 <=  20'h0cccd;
               12'b010001100110: data1 <=  20'h05095;
               12'b010001100111: data1 <=  20'h19094;
               12'b010001101000: data1 <=  20'h66126;
               12'b010001101001: data1 <=  20'h01cc9;
               12'b010001101010: data1 <=  20'h4f0e9;
               12'b010001101011: data1 <=  20'h849c3;
               12'b010001101100: data1 <=  20'h220c9;
               12'b010001101101: data1 <=  20'h21c8a;
               12'b010001101110: data1 <=  20'h280c9;
               12'b010001101111: data1 <=  20'h210c9;
               12'b010001110000: data1 <=  20'h5b144;
               12'b010001110001: data1 <=  20'h209ce;
               12'b010001110010: data1 <=  20'h35186;
               12'b010001110011: data1 <=  20'h2718c;
               12'b010001110100: data1 <=  20'h540ca;
               12'b010001110101: data1 <=  20'h3ee88;
               12'b010001110110: data1 <=  20'h55126;
               12'b010001110111: data1 <=  20'h024c9;
               12'b010001111000: data1 <=  20'h08cae;
               12'b010001111001: data1 <=  20'h19e06;
               12'b010001111010: data1 <=  20'h16d09;
               12'b010001111011: data1 <=  20'h530ca;
               12'b010001111100: data1 <=  20'h55126;
               12'b010001111101: data1 <=  20'h51526;
               12'b010001111110: data1 <=  20'h67526;
               12'b010001111111: data1 <=  20'h64926;
               12'b010010000000: data1 <=  20'h65643;
               12'b010010000001: data1 <=  20'h64643;
               12'b010010000010: data1 <=  20'h01643;
               12'b010010000011: data1 <=  20'h06a62;
               12'b010010000100: data1 <=  20'h100cb;
               12'b010010000101: data1 <=  20'h5ede6;
               12'b010010000110: data1 <=  20'h100cb;
               12'b010010000111: data1 <=  20'h0d8cb;
               12'b010010001000: data1 <=  20'h110c9;
               12'b010010001001: data1 <=  20'h0cec4;
               12'b010010001010: data1 <=  20'h00aac;
               12'b010010001011: data1 <=  20'h4b243;
               12'b010010001100: data1 <=  20'h0f8c9;
               12'b010010001101: data1 <=  20'h3f643;
               12'b010010001110: data1 <=  20'h16d09;
               12'b010010001111: data1 <=  20'h2ca43;
               12'b010010010000: data1 <=  20'h470c9;
               12'b010010010001: data1 <=  20'h344c9;
               12'b010010010010: data1 <=  20'h03c52;
               12'b010010010011: data1 <=  20'h01c52;
               12'b010010010100: data1 <=  20'h170e9;
               12'b010010010101: data1 <=  20'h71526;
               12'b010010010110: data1 <=  20'h716a3;
               12'b010010010111: data1 <=  20'h12ce9;
               12'b010010011000: data1 <=  20'h2c6c3;
               12'b010010011001: data1 <=  20'h12f10;
               12'b010010011010: data1 <=  20'h6d924;
               12'b010010011011: data1 <=  20'h20988;
               12'b010010011100: data1 <=  20'h26dc6;
               12'b010010011101: data1 <=  20'h655c6;
               12'b010010011110: data1 <=  20'h110c9;
               12'b010010011111: data1 <=  20'h0c8c9;
               12'b010010100000: data1 <=  20'h19e8a;
               12'b010010100001: data1 <=  20'h51d28;
               12'b010010100010: data1 <=  20'h06eaf;
               12'b010010100011: data1 <=  20'h4c5c8;
               12'b010010100100: data1 <=  20'h2d584;
               12'b010010100101: data1 <=  20'h20d26;
               12'b010010100110: data1 <=  20'h480c6;
               12'b010010100111: data1 <=  20'h460c6;
               12'b010010101000: data1 <=  20'h1aa42;
               12'b010010101001: data1 <=  20'h0c8cb;
               12'b010010101010: data1 <=  20'h048cf;
               12'b010010101011: data1 <=  20'h000cd;
               12'b010010101100: data1 <=  20'h030c9;
               12'b010010101101: data1 <=  20'h018c9;
               12'b010010101110: data1 <=  20'h0cb04;
               12'b010010101111: data1 <=  20'h52244;
               12'b010010110000: data1 <=  20'h2e144;
               12'b010010110001: data1 <=  20'h33583;
               12'b010010110010: data1 <=  20'h58a63;
               12'b010010110011: data1 <=  20'h02894;
               12'b010010110100: data1 <=  20'h5fd26;
               12'b010010110101: data1 <=  20'h38de4;
               12'b010010110110: data1 <=  20'h1b187;
               12'b010010110111: data1 <=  20'h3e8c9;
               12'b010010111000: data1 <=  20'h23cc9;
               12'b010010111001: data1 <=  20'h70a06;
               12'b010010111010: data1 <=  20'h72dc6;
               12'b010010111011: data1 <=  20'h7d684;
               12'b010010111100: data1 <=  20'h32a86;
               12'b010010111101: data1 <=  20'h33cc9;
               12'b010010111110: data1 <=  20'h21588;
               12'b010010111111: data1 <=  20'h20588;
               12'b010011000000: data1 <=  20'h280c9;
               12'b010011000001: data1 <=  20'h008d0;
               12'b010011000010: data1 <=  20'h1cccc;
               12'b010011000011: data1 <=  20'h19ccc;
               12'b010011000100: data1 <=  20'h4ed26;
               12'b010011000101: data1 <=  20'h011f6;
               12'b010011000110: data1 <=  20'h4ed26;
               12'b010011000111: data1 <=  20'h4b126;
               12'b010011001000: data1 <=  20'h61926;
               12'b010011001001: data1 <=  20'h5dd26;
               12'b010011001010: data1 <=  20'h0290a;
               12'b010011001011: data1 <=  20'h00490;
               12'b010011001100: data1 <=  20'h27546;
               12'b010011001101: data1 <=  20'h4d88a;
               12'b010011001110: data1 <=  20'h1b146;
               12'b010011001111: data1 <=  20'h8a642;
               12'b010011010000: data1 <=  20'h2d966;
               12'b010011010001: data1 <=  20'h0018a;
               12'b010011010010: data1 <=  20'h08d86;
               12'b010011010011: data1 <=  20'h65d24;
               12'b010011010100: data1 <=  20'h2d1f0;
               12'b010011010101: data1 <=  20'h3fd8d;
               12'b010011010110: data1 <=  20'h0e186;
               12'b010011010111: data1 <=  20'h39189;
               12'b010011011000: data1 <=  20'h10906;
               12'b010011011001: data1 <=  20'h0c906;
               12'b010011011010: data1 <=  20'h12f0b;
               12'b010011011011: data1 <=  20'h5150a;
               12'b010011011100: data1 <=  20'h5a08a;
               12'b010011011101: data1 <=  20'h0f095;
               12'b010011011110: data1 <=  20'h1a1e9;
               12'b010011011111: data1 <=  20'h06706;
               12'b010011100000: data1 <=  20'h27cb0;
               12'b010011100001: data1 <=  20'h84243;
               12'b010011100010: data1 <=  20'h20c6c;
               12'b010011100011: data1 <=  20'h28489;
               12'b010011100100: data1 <=  20'h26d28;
               12'b010011100101: data1 <=  20'h13e82;
               12'b010011100110: data1 <=  20'h3f243;
               12'b010011100111: data1 <=  20'h5f946;
               12'b010011101000: data1 <=  20'h19492;
               12'b010011101001: data1 <=  20'h034c9;
               12'b010011101010: data1 <=  20'h014c9;
               12'b010011101011: data1 <=  20'h02cc9;
               12'b010011101100: data1 <=  20'h2d526;
               12'b010011101101: data1 <=  20'h00e42;
               12'b010011101110: data1 <=  20'h3ea84;
               12'b010011101111: data1 <=  20'h0f08c;
               12'b010011110000: data1 <=  20'h20ccc;
               12'b010011110001: data1 <=  20'h01a56;
               12'b010011110010: data1 <=  20'h00256;
               12'b010011110011: data1 <=  20'h110cb;
               12'b010011110100: data1 <=  20'h0c8cb;
               12'b010011110101: data1 <=  20'h02cc9;
               12'b010011110110: data1 <=  20'h00283;
               12'b010011110111: data1 <=  20'h0d282;
               12'b010011111000: data1 <=  20'h3ee42;
               12'b010011111001: data1 <=  20'h304c9;
               12'b010011111010: data1 <=  20'h002c9;
               12'b010011111011: data1 <=  20'h170c9;
               12'b010011111100: data1 <=  20'h2bcc9;
               12'b010011111101: data1 <=  20'h25b06;
               12'b010011111110: data1 <=  20'h0c8ca;
               12'b010011111111: data1 <=  20'h280c9;
               12'b010100000000: data1 <=  20'h01cc9;
               12'b010100000001: data1 <=  20'h03cc9;
               12'b010100000010: data1 <=  20'h00cc9;
               12'b010100000011: data1 <=  20'h6e126;
               12'b010100000100: data1 <=  20'h6a643;
               12'b010100000101: data1 <=  20'h5b526;
               12'b010100000110: data1 <=  20'h5dee6;
               12'b010100000111: data1 <=  20'h5f243;
               12'b010100001000: data1 <=  20'h57926;
               12'b010100001001: data1 <=  20'h3450a;
               12'b010100001010: data1 <=  20'h2c9e6;
               12'b010100001011: data1 <=  20'h3450a;
               12'b010100001100: data1 <=  20'h014cc;
               12'b010100001101: data1 <=  20'h3450a;
               12'b010100001110: data1 <=  20'h214c9;
               12'b010100001111: data1 <=  20'h28092;
               12'b010100010000: data1 <=  20'h2d184;
               12'b010100010001: data1 <=  20'h3450a;
               12'b010100010010: data1 <=  20'h33d0a;
               12'b010100010011: data1 <=  20'h414ce;
               12'b010100010100: data1 <=  20'h218d3;
               12'b010100010101: data1 <=  20'h4c986;
               12'b010100010110: data1 <=  20'h38a46;
               12'b010100010111: data1 <=  20'h5b90a;
               12'b010100011000: data1 <=  20'h386c8;
               12'b010100011001: data1 <=  20'h72986;
               12'b010100011010: data1 <=  20'h25a92;
               12'b010100011011: data1 <=  20'h2668c;
               12'b010100011100: data1 <=  20'h64148;
               12'b010100011101: data1 <=  20'h65a43;
               12'b010100011110: data1 <=  20'h44e63;
               12'b010100011111: data1 <=  20'h290c9;
               12'b010100100000: data1 <=  20'h2c2c4;
               12'b010100100001: data1 <=  20'h28cec;
               12'b010100100010: data1 <=  20'h2cd69;
               12'b010100100011: data1 <=  20'h41948;
               12'b010100100100: data1 <=  20'h4b927;
               12'b010100100101: data1 <=  20'h5b8c9;
               12'b010100100110: data1 <=  20'h4bccc;
               12'b010100100111: data1 <=  20'h54cc6;
               12'b010100101000: data1 <=  20'h020c9;
               12'b010100101001: data1 <=  20'h088d7;
               12'b010100101010: data1 <=  20'h64126;
               12'b010100101011: data1 <=  20'h6b643;
               12'b010100101100: data1 <=  20'h0ddae;
               12'b010100101101: data1 <=  20'h03d0c;
               12'b010100101110: data1 <=  20'h0010c;
               12'b010100101111: data1 <=  20'h0e907;
               12'b010100110000: data1 <=  20'h068c9;
               12'b010100110001: data1 <=  20'h358cc;
               12'b010100110010: data1 <=  20'h330cc;
               12'b010100110011: data1 <=  20'h234af;
               12'b010100110100: data1 <=  20'h200af;
               12'b010100110101: data1 <=  20'h1d8c9;
               12'b010100110110: data1 <=  20'h2c0cf;
               12'b010100110111: data1 <=  20'h60988;
               12'b010100111000: data1 <=  20'h0cb04;
               12'b010100111001: data1 <=  20'h0a053;
               12'b010100111010: data1 <=  20'h08053;
               12'b010100111011: data1 <=  20'h0bc54;
               12'b010100111100: data1 <=  20'h06454;
               12'b010100111101: data1 <=  20'h494cc;
               12'b010100111110: data1 <=  20'h44ccc;
               12'b010100111111: data1 <=  20'h2664e;
               12'b010101000000: data1 <=  20'h400e8;
               12'b010101000001: data1 <=  20'h3a18c;
               12'b010101000010: data1 <=  20'h71245;
               12'b010101000011: data1 <=  20'h84683;
               12'b010101000100: data1 <=  20'h4d4cc;
               12'b010101000101: data1 <=  20'h26a43;
               12'b010101000110: data1 <=  20'h26643;
               12'b010101000111: data1 <=  20'h1d8c9;
               12'b010101001000: data1 <=  20'h4b926;
               12'b010101001001: data1 <=  20'h58a44;
               12'b010101001010: data1 <=  20'h2d8ce;
               12'b010101001011: data1 <=  20'h53186;
               12'b010101001100: data1 <=  20'h2d589;
               12'b010101001101: data1 <=  20'h4e0c6;
               12'b010101001110: data1 <=  20'h0c88a;
               12'b010101001111: data1 <=  20'h02126;
               12'b010101010000: data1 <=  20'h38d86;
               12'b010101010001: data1 <=  20'h41cc9;
               12'b010101010010: data1 <=  20'h3fcc9;
               12'b010101010011: data1 <=  20'h60126;
               12'b010101010100: data1 <=  20'h65586;
               12'b010101010101: data1 <=  20'h0d683;
               12'b010101010110: data1 <=  20'h1fd86;
               12'b010101010111: data1 <=  20'h02c78;
               12'b010101011000: data1 <=  20'h64de4;
               12'b010101011001: data1 <=  20'h4d4cc;
               12'b010101011010: data1 <=  20'h5e188;
               12'b010101011011: data1 <=  20'h4250e;
               12'b010101011100: data1 <=  20'h3890e;
               12'b010101011101: data1 <=  20'h4712a;
               12'b010101011110: data1 <=  20'h2d586;
               12'b010101011111: data1 <=  20'h604c9;
               12'b010101100000: data1 <=  20'h33d27;
               12'b010101100001: data1 <=  20'h1b90a;
               12'b010101100010: data1 <=  20'h268c9;
               12'b010101100011: data1 <=  20'h25b0c;
               12'b010101100100: data1 <=  20'h2c8ce;
               12'b010101100101: data1 <=  20'h36ca8;
               12'b010101100110: data1 <=  20'h320a8;
               12'b010101100111: data1 <=  20'h170c6;
               12'b010101101000: data1 <=  20'h130c6;
               12'b010101101001: data1 <=  20'h110c9;
               12'b010101101010: data1 <=  20'h0c8c9;
               12'b010101101011: data1 <=  20'h13a46;
               12'b010101101100: data1 <=  20'h13526;
               12'b010101101101: data1 <=  20'h15148;
               12'b010101101110: data1 <=  20'h14148;
               12'b010101101111: data1 <=  20'h474cc;
               12'b010101110000: data1 <=  20'h46ccb;
               12'b010101110001: data1 <=  20'h33d44;
               12'b010101110010: data1 <=  20'h27cc7;
               12'b010101110011: data1 <=  20'h71e43;
               12'b010101110100: data1 <=  20'h1b0c9;
               12'b010101110101: data1 <=  20'h08527;
               12'b010101110110: data1 <=  20'h464c6;
               12'b010101110111: data1 <=  20'h4e88b;
               12'b010101111000: data1 <=  20'h4c88b;
               12'b010101111001: data1 <=  20'h02192;
               12'b010101111010: data1 <=  20'h4b945;
               12'b010101111011: data1 <=  20'h7dac3;
               12'b010101111100: data1 <=  20'h19054;
               12'b010101111101: data1 <=  20'h0cb04;
               12'b010101111110: data1 <=  20'h33d44;
               12'b010101111111: data1 <=  20'h2d50a;
               12'b010110000000: data1 <=  20'h038ce;
               12'b010110000001: data1 <=  20'h45ca8;
               12'b010110000010: data1 <=  20'h00a89;
               12'b010110000011: data1 <=  20'h2d588;
               12'b010110000100: data1 <=  20'h6c8c6;
               12'b010110000101: data1 <=  20'h40544;
               12'b010110000110: data1 <=  20'h20d89;
               12'b010110000111: data1 <=  20'h460c8;
               12'b010110001000: data1 <=  20'h1d891;
               12'b010110001001: data1 <=  20'h000c6;
               12'b010110001010: data1 <=  20'h1d891;
               12'b010110001011: data1 <=  20'h19891;
               12'b010110001100: data1 <=  20'h71e63;
               12'b010110001101: data1 <=  20'h02c52;
               12'b010110001110: data1 <=  20'h1cc52;
               12'b010110001111: data1 <=  20'h1ac52;
               12'b010110010000: data1 <=  20'h46948;
               12'b010110010001: data1 <=  20'h28089;
               12'b010110010010: data1 <=  20'h028c9;
               12'b010110010011: data1 <=  20'h38e08;
               12'b010110010100: data1 <=  20'h614c9;
               12'b010110010101: data1 <=  20'h2dcc9;
               12'b010110010110: data1 <=  20'h614c9;
               12'b010110010111: data1 <=  20'h4bd86;
               12'b010110011000: data1 <=  20'h4e926;
               12'b010110011001: data1 <=  20'h4b526;
               12'b010110011010: data1 <=  20'h2ca43;
               12'b010110011011: data1 <=  20'h2c2c6;
               12'b010110011100: data1 <=  20'h1d8c6;
               12'b010110011101: data1 <=  20'h190c6;
               12'b010110011110: data1 <=  20'h46206;
               12'b010110011111: data1 <=  20'h65924;
               12'b010110100000: data1 <=  20'h614c9;
               12'b010110100001: data1 <=  20'h5ecc9;
               12'b010110100010: data1 <=  20'h0a0d7;
               12'b010110100011: data1 <=  20'h83703;
               12'b010110100100: data1 <=  20'h7d304;
               12'b010110100101: data1 <=  20'h070d7;
               12'b010110100110: data1 <=  20'h6b243;
               12'b010110100111: data1 <=  20'h64243;
               12'b010110101000: data1 <=  20'h646c4;
               12'b010110101001: data1 <=  20'h64126;
               12'b010110101010: data1 <=  20'h3f2a3;
               12'b010110101011: data1 <=  20'h71186;
               12'b010110101100: data1 <=  20'h1f704;
               12'b010110101101: data1 <=  20'h0f08f;
               12'b010110101110: data1 <=  20'h2e4cc;
               12'b010110101111: data1 <=  20'h270c9;
               12'b010110110000: data1 <=  20'h02cc9;
               12'b010110110001: data1 <=  20'h2e0c9;
               12'b010110110010: data1 <=  20'h06e83;
               12'b010110110011: data1 <=  20'h70d86;
               12'b010110110100: data1 <=  20'h0fc8d;
               12'b010110110101: data1 <=  20'h2d584;
               12'b010110110110: data1 <=  20'h08c8d;
               12'b010110110111: data1 <=  20'h01872;
               12'b010110111000: data1 <=  20'h16545;
               12'b010110111001: data1 <=  20'h5f588;
               12'b010110111010: data1 <=  20'h40cc9;
               12'b010110111011: data1 <=  20'h14c89;
               12'b010110111100: data1 <=  20'h044ce;
               12'b010110111101: data1 <=  20'h004ce;
               12'b010110111110: data1 <=  20'h038d0;
               12'b010110111111: data1 <=  20'h1ac8a;
               12'b010111000000: data1 <=  20'h6b246;
               12'b010111000001: data1 <=  20'h7d6c4;
               12'b010111000010: data1 <=  20'h16545;
               12'b010111000011: data1 <=  20'h12d45;
               12'b010111000100: data1 <=  20'h28990;
               12'b010111000101: data1 <=  20'h25990;
               12'b010111000110: data1 <=  20'h3acaf;
               12'b010111000111: data1 <=  20'h70ea2;
               12'b010111001000: data1 <=  20'h03d26;
               12'b010111001001: data1 <=  20'h07d84;
               12'b010111001010: data1 <=  20'h0198c;
               12'b010111001011: data1 <=  20'h4090c;
               12'b010111001100: data1 <=  20'h67948;
               12'b010111001101: data1 <=  20'h64148;
               12'b010111001110: data1 <=  20'h4d985;
               12'b010111001111: data1 <=  20'h65948;
               12'b010111010000: data1 <=  20'h27586;
               12'b010111010001: data1 <=  20'h27c92;
               12'b010111010010: data1 <=  20'h3acce;
               12'b010111010011: data1 <=  20'h3a4ce;
               12'b010111010100: data1 <=  20'h1ad6c;
               12'b010111010101: data1 <=  20'h330d0;
               12'b010111010110: data1 <=  20'h17095;
               12'b010111010111: data1 <=  20'h13895;
               12'b010111011000: data1 <=  20'h08d12;
               12'b010111011001: data1 <=  20'h1fe08;
               12'b010111011010: data1 <=  20'h2664c;
               12'b010111011011: data1 <=  20'h3fa0c;
               12'b010111011100: data1 <=  20'h1cd14;
               12'b010111011101: data1 <=  20'h0e526;
               12'b010111011110: data1 <=  20'h1cd14;
               12'b010111011111: data1 <=  20'h19514;
               12'b010111100000: data1 <=  20'h34d0e;
               12'b010111100001: data1 <=  20'h3350e;
               12'b010111100010: data1 <=  20'h53ca8;
               12'b010111100011: data1 <=  20'h524e9;
               12'b010111100100: data1 <=  20'h5170a;
               12'b010111100101: data1 <=  20'h0d90b;
               12'b010111100110: data1 <=  20'h0f110;
               12'b010111100111: data1 <=  20'h0cb06;
               12'b010111101000: data1 <=  20'h01989;
               12'b010111101001: data1 <=  20'h0cd8c;
               12'b010111101010: data1 <=  20'h23cc9;
               12'b010111101011: data1 <=  20'h13d0a;
               12'b010111101100: data1 <=  20'h84e43;
               12'b010111101101: data1 <=  20'h3ee42;
               12'b010111101110: data1 <=  20'h3eec3;
               12'b010111101111: data1 <=  20'h32989;
               12'b010111110000: data1 <=  20'h35186;
               12'b010111110001: data1 <=  20'h32186;
               12'b010111110010: data1 <=  20'h604c9;
               12'b010111110011: data1 <=  20'h53126;
               12'b010111110100: data1 <=  20'h344ec;
               12'b010111110101: data1 <=  20'h52526;
               12'b010111110110: data1 <=  20'h5f644;
               12'b010111110111: data1 <=  20'h1a490;
               12'b010111111000: data1 <=  20'h604c9;
               12'b010111111001: data1 <=  20'h5fcc9;
               12'b010111111010: data1 <=  20'h4718a;
               12'b010111111011: data1 <=  20'h265c6;
               12'b010111111100: data1 <=  20'h0da28;
               12'b010111111101: data1 <=  20'h0e195;
               12'b010111111110: data1 <=  20'h08529;
               12'b010111111111: data1 <=  20'h2bf03;
               12'b011000000000: data1 <=  20'h2852a;
               12'b011000000001: data1 <=  20'h45643;
               12'b011000000010: data1 <=  20'h66124;
               12'b011000000011: data1 <=  20'h00126;
               12'b011000000100: data1 <=  20'h44f06;
               12'b011000000101: data1 <=  20'h38e86;
               12'b011000000110: data1 <=  20'h2060c;
               12'b011000000111: data1 <=  20'h0f08f;
               12'b011000001000: data1 <=  20'h14944;
               12'b011000001001: data1 <=  20'h600c8;
               12'b011000001010: data1 <=  20'h044ea;
               12'b011000001011: data1 <=  20'h000ea;
               12'b011000001100: data1 <=  20'h0a4cc;
               12'b011000001101: data1 <=  20'h00668;
               12'b011000001110: data1 <=  20'h0f924;
               12'b011000001111: data1 <=  20'h0d524;
               12'b011000010000: data1 <=  20'h0f946;
               12'b011000010001: data1 <=  20'h19e42;
               12'b011000010010: data1 <=  20'h09489;
               12'b011000010011: data1 <=  20'h08489;
               12'b011000010100: data1 <=  20'h21d0a;
               12'b011000010101: data1 <=  20'h1a98d;
               12'b011000010110: data1 <=  20'h228c6;
               12'b011000010111: data1 <=  20'h1f983;
               12'b011000011000: data1 <=  20'h21146;
               12'b011000011001: data1 <=  20'h00aa5;
               12'b011000011010: data1 <=  20'h32129;
               12'b011000011011: data1 <=  20'h27cc9;
               12'b011000011100: data1 <=  20'h12cc7;
               12'b011000011101: data1 <=  20'h72d86;
               12'b011000011110: data1 <=  20'h32a86;
               12'b011000011111: data1 <=  20'h0fd44;
               12'b011000100000: data1 <=  20'h204b2;
               12'b011000100001: data1 <=  20'h1e089;
               12'b011000100010: data1 <=  20'h2790e;
               12'b011000100011: data1 <=  20'h06706;
               12'b011000100100: data1 <=  20'h19089;
               12'b011000100101: data1 <=  20'h26643;
               12'b011000100110: data1 <=  20'h6b206;
               12'b011000100111: data1 <=  20'h28cc9;
               12'b011000101000: data1 <=  20'h26dc6;
               12'b011000101001: data1 <=  20'h2290a;
               12'b011000101010: data1 <=  20'h0d283;
               12'b011000101011: data1 <=  20'h0ed26;
               12'b011000101100: data1 <=  20'h278c9;
               12'b011000101101: data1 <=  20'h15c8b;
               12'b011000101110: data1 <=  20'h14c8b;
               12'b011000101111: data1 <=  20'h14d0a;
               12'b011000110000: data1 <=  20'h09052;
               12'b011000110001: data1 <=  20'h0ed26;
               12'b011000110010: data1 <=  20'h0ca63;
               12'b011000110011: data1 <=  20'h59d26;
               12'b011000110100: data1 <=  20'h32645;
               12'b011000110101: data1 <=  20'h030c9;
               12'b011000110110: data1 <=  20'h018c9;
               12'b011000110111: data1 <=  20'h28c8f;
               12'b011000111000: data1 <=  20'h1fa43;
               12'b011000111001: data1 <=  20'h2e1c6;
               12'b011000111010: data1 <=  20'h64a43;
               12'b011000111011: data1 <=  20'h6e126;
               12'b011000111100: data1 <=  20'h32186;
               12'b011000111101: data1 <=  20'h538e8;
               12'b011000111110: data1 <=  20'h6ae83;
               12'b011000111111: data1 <=  20'h6e126;
               12'b011001000000: data1 <=  20'h011e4;
               12'b011001000001: data1 <=  20'h10cc6;
               12'b011001000010: data1 <=  20'h12cc9;
               12'b011001000011: data1 <=  20'h6e126;
               12'b011001000100: data1 <=  20'h6a526;
               12'b011001000101: data1 <=  20'h72d86;
               12'b011001000110: data1 <=  20'h5e8c9;
               12'b011001000111: data1 <=  20'h5550a;
               12'b011001001000: data1 <=  20'h57b04;
               12'b011001001001: data1 <=  20'h73cc6;
               12'b011001001010: data1 <=  20'h5150a;
               12'b011001001011: data1 <=  20'h57b06;
               12'b011001001100: data1 <=  20'h0dd88;
               12'b011001001101: data1 <=  20'h3a526;
               12'b011001001110: data1 <=  20'h13e04;
               12'b011001001111: data1 <=  20'h0f08a;
               12'b011001010000: data1 <=  20'h1b0a8;
               12'b011001010001: data1 <=  20'h2212c;
               12'b011001010010: data1 <=  20'h2052c;
               12'b011001010011: data1 <=  20'h290c9;
               12'b011001010100: data1 <=  20'h19a8c;
               12'b011001010101: data1 <=  20'h1a230;
               12'b011001010110: data1 <=  20'h2dce6;
               12'b011001010111: data1 <=  20'h38ae2;
               12'b011001011000: data1 <=  20'h01cc9;
               12'b011001011001: data1 <=  20'h16089;
               12'b011001011010: data1 <=  20'h084cd;
               12'b011001011011: data1 <=  20'h8aa42;
               12'b011001011100: data1 <=  20'h3f526;
               12'b011001011101: data1 <=  20'h03858;
               12'b011001011110: data1 <=  20'h02058;
               12'b011001011111: data1 <=  20'h0d64a;
               12'b011001100000: data1 <=  20'h525e6;
               12'b011001100001: data1 <=  20'h84243;
               12'b011001100010: data1 <=  20'h0888b;
               12'b011001100011: data1 <=  20'h2e144;
               12'b011001100100: data1 <=  20'h01d52;
               12'b011001100101: data1 <=  20'h094d0;
               12'b011001100110: data1 <=  20'h07cd0;
               12'b011001100111: data1 <=  20'h110c6;
               12'b011001101000: data1 <=  20'h20242;
               12'b011001101001: data1 <=  20'h110c6;
               12'b011001101010: data1 <=  20'h0c8c6;
               12'b011001101011: data1 <=  20'h48166;
               12'b011001101100: data1 <=  20'h2d144;
               12'b011001101101: data1 <=  20'h3b147;
               12'b011001101110: data1 <=  20'h39147;
               12'b011001101111: data1 <=  20'h1d0c6;
               12'b011001110000: data1 <=  20'h26d48;
               12'b011001110001: data1 <=  20'h85203;
               12'b011001110010: data1 <=  20'h83a03;
               12'b011001110011: data1 <=  20'h1fece;
               12'b011001110100: data1 <=  20'h3f50a;
               12'b011001110101: data1 <=  20'h044cc;
               12'b011001110110: data1 <=  20'h0dcd2;
               12'b011001110111: data1 <=  20'h034c9;
               12'b011001111000: data1 <=  20'h4b0e9;
               12'b011001111001: data1 <=  20'h5510a;
               12'b011001111010: data1 <=  20'h004cc;
               12'b011001111011: data1 <=  20'h0946c;
               12'b011001111100: data1 <=  20'h5190a;
               12'b011001111101: data1 <=  20'h84262;
               12'b011001111110: data1 <=  20'h1448d;
               12'b011001111111: data1 <=  20'h3fe43;
               12'b011010000000: data1 <=  20'h150ac;
               12'b011010000001: data1 <=  20'h0f48f;
               12'b011010000010: data1 <=  20'h07604;
               12'b011010000011: data1 <=  20'h01a43;
               12'b011010000100: data1 <=  20'h07948;
               12'b011010000101: data1 <=  20'h73586;
               12'b011010000110: data1 <=  20'h5f183;
               12'b011010000111: data1 <=  20'h3eec4;
               12'b011010001000: data1 <=  20'h3a126;
               12'b011010001001: data1 <=  20'h46585;
               12'b011010001010: data1 <=  20'h2d547;
               12'b011010001011: data1 <=  20'h0f50a;
               12'b011010001100: data1 <=  20'h0dd0a;
               12'b011010001101: data1 <=  20'h1aa46;
               12'b011010001110: data1 <=  20'h1f549;
               12'b011010001111: data1 <=  20'h2c6a6;
               12'b011010010000: data1 <=  20'h192d0;
               12'b011010010001: data1 <=  20'h024d6;
               12'b011010010010: data1 <=  20'h0886c;
               12'b011010010011: data1 <=  20'h03192;
               12'b011010010100: data1 <=  20'h00192;
               12'b011010010101: data1 <=  20'h06ac4;
               12'b011010010110: data1 <=  20'h00e44;
               12'b011010010111: data1 <=  20'h1fec6;
               12'b011010011000: data1 <=  20'h014c9;
               12'b011010011001: data1 <=  20'h5a0c9;
               12'b011010011010: data1 <=  20'h598c9;
               12'b011010011011: data1 <=  20'h71e43;
               12'b011010011100: data1 <=  20'h018cd;
               12'b011010011101: data1 <=  20'h1ad84;
               12'b011010011110: data1 <=  20'h0dd86;
               12'b011010011111: data1 <=  20'h07643;
               12'b011010100000: data1 <=  20'h320cc;
               12'b011010100001: data1 <=  20'h600c9;
               12'b011010100010: data1 <=  20'h40ccd;
               12'b011010100011: data1 <=  20'h6be42;
               12'b011010100100: data1 <=  20'h1b4c9;
               12'b011010100101: data1 <=  20'h028c9;
               12'b011010100110: data1 <=  20'h26d48;
               12'b011010100111: data1 <=  20'h3bca8;
               12'b011010101000: data1 <=  20'h398a8;
               12'b011010101001: data1 <=  20'h48526;
               12'b011010101010: data1 <=  20'h0caef;
               12'b011010101011: data1 <=  20'h0410c;
               12'b011010101100: data1 <=  20'h5ecc9;
               12'b011010101101: data1 <=  20'h72924;
               12'b011010101110: data1 <=  20'h6a643;
               12'b011010101111: data1 <=  20'h48166;
               12'b011010110000: data1 <=  20'h44d66;
               12'b011010110001: data1 <=  20'h38706;
               12'b011010110010: data1 <=  20'h65908;
               12'b011010110011: data1 <=  20'h669c6;
               12'b011010110100: data1 <=  20'h06aa3;
               12'b011010110101: data1 <=  20'h0cb03;
               12'b011010110110: data1 <=  20'h5e505;
               12'b011010110111: data1 <=  20'h456a3;
               12'b011010111000: data1 <=  20'h70d86;
               12'b011010111001: data1 <=  20'h5a08a;
               12'b011010111010: data1 <=  20'h2d88a;
               12'b011010111011: data1 <=  20'h344cc;
               12'b011010111100: data1 <=  20'h08126;
               12'b011010111101: data1 <=  20'h58662;
               12'b011010111110: data1 <=  20'h2d94a;
               12'b011010111111: data1 <=  20'h4be4c;
               12'b011011000000: data1 <=  20'h020cc;
               12'b011011000001: data1 <=  20'h00e29;
               12'b011011000010: data1 <=  20'h0198b;
               12'b011011000011: data1 <=  20'h004cd;
               12'b011011000100: data1 <=  20'h33606;
               12'b011011000101: data1 <=  20'h340ac;
               12'b011011000110: data1 <=  20'h84243;
               12'b011011000111: data1 <=  20'h000c6;
               12'b011011001000: data1 <=  20'h00a83;
               12'b011011001001: data1 <=  20'h269ea;
               12'b011011001010: data1 <=  20'h27cc9;
               12'b011011001011: data1 <=  20'h024c9;
               12'b011011001100: data1 <=  20'h038c9;
               12'b011011001101: data1 <=  20'h65d26;
               12'b011011001110: data1 <=  20'h038c9;
               12'b011011001111: data1 <=  20'h010c9;
               12'b011011010000: data1 <=  20'h0a8d0;
               12'b011011010001: data1 <=  20'h068d0;
               12'b011011010010: data1 <=  20'h54cc9;
               12'b011011010011: data1 <=  20'h000c9;
               12'b011011010100: data1 <=  20'h218c6;
               12'b011011010101: data1 <=  20'h3f526;
               12'b011011010110: data1 <=  20'h2f470;
               12'b011011010111: data1 <=  20'h3f9cc;
               12'b011011011000: data1 <=  20'h27586;
               12'b011011011001: data1 <=  20'h0e494;
               12'b011011011010: data1 <=  20'h54cc9;
               12'b011011011011: data1 <=  20'h28089;
               12'b011011011100: data1 <=  20'h54cc9;
               12'b011011011101: data1 <=  20'h7e5c4;
               12'b011011011110: data1 <=  20'h1a20c;
               12'b011011011111: data1 <=  20'h27cc9;
               12'b011011100000: data1 <=  20'h00ea4;
               12'b011011100001: data1 <=  20'h524c9;
               12'b011011100010: data1 <=  20'h680a8;
               12'b011011100011: data1 <=  20'h01210;
               12'b011011100100: data1 <=  20'h271c6;
               12'b011011100101: data1 <=  20'h21c8f;
               12'b011011100110: data1 <=  20'h60188;
               12'b011011100111: data1 <=  20'h2d584;
               12'b011011101000: data1 <=  20'h26dc6;
               12'b011011101001: data1 <=  20'h2664a;
               12'b011011101010: data1 <=  20'h01a55;
               12'b011011101011: data1 <=  20'h00315;
               12'b011011101100: data1 <=  20'h72243;
               12'b011011101101: data1 <=  20'h5dd26;
               12'b011011101110: data1 <=  20'h13e62;
               12'b011011101111: data1 <=  20'h12f02;
               12'b011011110000: data1 <=  20'h5b524;
               12'b011011110001: data1 <=  20'h57924;
               12'b011011110010: data1 <=  20'h5f642;
               12'b011011110011: data1 <=  20'h6b243;
               12'b011011110100: data1 <=  20'h03077;
               12'b011011110101: data1 <=  20'h01906;
               12'b011011110110: data1 <=  20'h65a43;
               12'b011011110111: data1 <=  20'h02477;
               12'b011011111000: data1 <=  20'h2e48a;
               12'b011011111001: data1 <=  20'h33d4c;
               12'b011011111010: data1 <=  20'h3bcce;
               12'b011011111011: data1 <=  20'h00949;
               12'b011011111100: data1 <=  20'h090ac;
               12'b011011111101: data1 <=  20'h1958a;
               12'b011011111110: data1 <=  20'h0a124;
               12'b011011111111: data1 <=  20'h0cd0a;
               12'b011100000000: data1 <=  20'h08cac;
               12'b011100000001: data1 <=  20'h011d8;
               12'b011100000010: data1 <=  20'h6c144;
               12'b011100000011: data1 <=  20'h5a08a;
               12'b011100000100: data1 <=  20'h610c9;
               12'b011100000101: data1 <=  20'h84243;
               12'b011100000110: data1 <=  20'h610c9;
               12'b011100000111: data1 <=  20'h5f0c9;
               12'b011100001000: data1 <=  20'h28092;
               12'b011100001001: data1 <=  20'h148cb;
               12'b011100001010: data1 <=  20'h0a124;
               12'b011100001011: data1 <=  20'h1a5c8;
               12'b011100001100: data1 <=  20'h085e9;
               12'b011100001101: data1 <=  20'h0e50a;
               12'b011100001110: data1 <=  20'h0f8cc;
               12'b011100001111: data1 <=  20'h0e0cc;
               12'b011100010000: data1 <=  20'h2d984;
               12'b011100010001: data1 <=  20'h1458a;
               12'b011100010010: data1 <=  20'h26e06;
               12'b011100010011: data1 <=  20'h07249;
               12'b011100010100: data1 <=  20'h32e45;
               12'b011100010101: data1 <=  20'h00316;
               12'b011100010110: data1 <=  20'h67926;
               12'b011100010111: data1 <=  20'h64308;
               12'b011100011000: data1 <=  20'h772c4;
               12'b011100011001: data1 <=  20'h64526;
               12'b011100011010: data1 <=  20'h33d44;
               12'b011100011011: data1 <=  20'h600c9;
               12'b011100011100: data1 <=  20'h73186;
               12'b011100011101: data1 <=  20'h71186;
               12'b011100011110: data1 <=  20'h14e09;
               12'b011100011111: data1 <=  20'h1f546;
               12'b011100100000: data1 <=  20'h20a43;
               12'b011100100001: data1 <=  20'h26126;
               12'b011100100010: data1 <=  20'h10149;
               12'b011100100011: data1 <=  20'h26643;
               12'b011100100100: data1 <=  20'h0ede6;
               12'b011100100101: data1 <=  20'h331e6;
               12'b011100100110: data1 <=  20'h1f704;
               12'b011100100111: data1 <=  20'h33ccc;
               12'b011100101000: data1 <=  20'h02cc9;
               12'b011100101001: data1 <=  20'h4b0cc;
               12'b011100101010: data1 <=  20'h4e946;
               12'b011100101011: data1 <=  20'h2c649;
               12'b011100101100: data1 <=  20'h5a549;
               12'b011100101101: data1 <=  20'h27548;
               12'b011100101110: data1 <=  20'h271c6;
               12'b011100101111: data1 <=  20'h52527;
               12'b011100110000: data1 <=  20'h420cc;
               12'b011100110001: data1 <=  20'h3f8cc;
               12'b011100110010: data1 <=  20'h3b906;
               12'b011100110011: data1 <=  20'h14c8e;
               12'b011100110100: data1 <=  20'h04472;
               12'b011100110101: data1 <=  20'h4c20c;
               12'b011100110110: data1 <=  20'h03cce;
               12'b011100110111: data1 <=  20'h00cce;
               12'b011100111000: data1 <=  20'h0f994;
               12'b011100111001: data1 <=  20'h0c994;
               12'b011100111010: data1 <=  20'h040d1;
               12'b011100111011: data1 <=  20'h008d1;
               12'b011100111100: data1 <=  20'h29526;
               12'b011100111101: data1 <=  20'h25926;
               12'b011100111110: data1 <=  20'h0accd;
               12'b011100111111: data1 <=  20'h064cd;
               12'b011101000000: data1 <=  20'h04089;
               12'b011101000001: data1 <=  20'h3fd87;
               12'b011101000010: data1 <=  20'h3b586;
               12'b011101000011: data1 <=  20'h38586;
               12'b011101000100: data1 <=  20'h2d1c9;
               12'b011101000101: data1 <=  20'h5de83;
               12'b011101000110: data1 <=  20'h4090a;
               12'b011101000111: data1 <=  20'h1a5a9;
               12'b011101001000: data1 <=  20'h0f0d2;
               12'b011101001001: data1 <=  20'h018c9;
               12'b011101001010: data1 <=  20'h39d84;
               12'b011101001011: data1 <=  20'h0d5ec;
               12'b011101001100: data1 <=  20'h03185;
               12'b011101001101: data1 <=  20'h5de43;
               12'b011101001110: data1 <=  20'h57b05;
               12'b011101001111: data1 <=  20'h07872;
               12'b011101010000: data1 <=  20'h0288e;
               12'b011101010001: data1 <=  20'h15089;
               12'b011101010010: data1 <=  20'h0e986;
               12'b011101010011: data1 <=  20'h19224;
               12'b011101010100: data1 <=  20'h680a8;
               12'b011101010101: data1 <=  20'h64ca8;
               12'b011101010110: data1 <=  20'h72242;
               12'b011101010111: data1 <=  20'h00185;
               12'b011101011000: data1 <=  20'h164cc;
               12'b011101011001: data1 <=  20'h4b0cc;
               12'b011101011010: data1 <=  20'h136a3;
               12'b011101011011: data1 <=  20'h13ccc;
               12'b011101011100: data1 <=  20'h35186;
               12'b011101011101: data1 <=  20'h5de09;
               12'b011101011110: data1 <=  20'h52e45;
               12'b011101011111: data1 <=  20'h25de6;
               12'b011101100000: data1 <=  20'h3b126;
               12'b011101100001: data1 <=  20'h00deb;
               12'b011101100010: data1 <=  20'h16872;
               12'b011101100011: data1 <=  20'h14472;
               12'b011101100100: data1 <=  20'h21948;
               12'b011101100101: data1 <=  20'h1a208;
               12'b011101100110: data1 <=  20'h2d983;
               12'b011101100111: data1 <=  20'h0152d;
               12'b011101101000: data1 <=  20'h02cc9;
               12'b011101101001: data1 <=  20'h01cc9;
               12'b011101101010: data1 <=  20'h08549;
               12'b011101101011: data1 <=  20'h0ca42;
               12'b011101101100: data1 <=  20'h53dc6;
               12'b011101101101: data1 <=  20'h515c6;
               12'b011101101110: data1 <=  20'h11875;
               12'b011101101111: data1 <=  20'h384ac;
               12'b011101110000: data1 <=  20'h28986;
               12'b011101110001: data1 <=  20'h32683;
               12'b011101110010: data1 <=  20'h2d263;
               12'b011101110011: data1 <=  20'h4b526;
               12'b011101110100: data1 <=  20'h401cc;
               12'b011101110101: data1 <=  20'h26dd2;
               12'b011101110110: data1 <=  20'h4dd27;
               12'b011101110111: data1 <=  20'h5e244;
               12'b011101111000: data1 <=  20'h5a4c9;
               12'b011101111001: data1 <=  20'h32244;
               12'b011101111010: data1 <=  20'h3f686;
               12'b011101111011: data1 <=  20'h3ee86;
               12'b011101111100: data1 <=  20'h38702;
               12'b011101111101: data1 <=  20'h4b688;
               12'b011101111110: data1 <=  20'h4dd27;
               12'b011101111111: data1 <=  20'h4c127;
               12'b011110000000: data1 <=  20'h4e105;
               12'b011110000001: data1 <=  20'h4c105;
               12'b011110000010: data1 <=  20'h41c8a;
               12'b011110000011: data1 <=  20'h5e282;
               12'b011110000100: data1 <=  20'h40cc6;
               12'b011110000101: data1 <=  20'h066a3;
               12'b011110000110: data1 <=  20'h1a9a9;
               12'b011110000111: data1 <=  20'h20d85;
               12'b011110001000: data1 <=  20'h41146;
               12'b011110001001: data1 <=  20'h4c8a8;
               12'b011110001010: data1 <=  20'h034c9;
               12'b011110001011: data1 <=  20'h3f246;
               12'b011110001100: data1 <=  20'h0f524;
               12'b011110001101: data1 <=  20'h7d6a3;
               12'b011110001110: data1 <=  20'h3eec2;
               12'b011110001111: data1 <=  20'h6a643;
               12'b011110010000: data1 <=  20'h034c9;
               12'b011110010001: data1 <=  20'h014c9;
               12'b011110010010: data1 <=  20'h110d4;
               12'b011110010011: data1 <=  20'h0c8d4;
               12'b011110010100: data1 <=  20'h2e8ce;
               12'b011110010101: data1 <=  20'h06489;
               12'b011110010110: data1 <=  20'h5a924;
               12'b011110010111: data1 <=  20'h51924;
               12'b011110011000: data1 <=  20'h275e6;
               12'b011110011001: data1 <=  20'h0e872;
               12'b011110011010: data1 <=  20'h27186;
               12'b011110011011: data1 <=  20'h77684;
               12'b011110011100: data1 <=  20'h614c9;
               12'b011110011101: data1 <=  20'h2024e;
               12'b011110011110: data1 <=  20'h29492;
               12'b011110011111: data1 <=  20'h26c92;
               12'b011110100000: data1 <=  20'h02cc9;
               12'b011110100001: data1 <=  20'h01cc9;
               12'b011110100010: data1 <=  20'h220c9;
               12'b011110100011: data1 <=  20'h218c6;
               12'b011110100100: data1 <=  20'h07606;
               12'b011110100101: data1 <=  20'h538cb;
               12'b011110100110: data1 <=  20'h0a8cc;
               12'b011110100111: data1 <=  20'h6aa43;
               12'b011110101000: data1 <=  20'h53148;
               12'b011110101001: data1 <=  20'h72146;
               12'b011110101010: data1 <=  20'h59d24;
               12'b011110101011: data1 <=  20'h068cc;
               12'b011110101100: data1 <=  20'h1dcac;
               12'b011110101101: data1 <=  20'h00108;
               12'b011110101110: data1 <=  20'h20263;
               12'b011110101111: data1 <=  20'h1f986;
               12'b011110110000: data1 <=  20'h06ea8;
               12'b011110110001: data1 <=  20'h07608;
               12'b011110110010: data1 <=  20'h01a43;
               12'b011110110011: data1 <=  20'h1a14e;
               12'b011110110100: data1 <=  20'h2948a;
               12'b011110110101: data1 <=  20'h71643;
               12'b011110110110: data1 <=  20'h72986;
               12'b011110110111: data1 <=  20'h5e8c9;
               12'b011110111000: data1 <=  20'h2f8c8;
               12'b011110111001: data1 <=  20'h2c8c8;
               12'b011110111010: data1 <=  20'h39a46;
               12'b011110111011: data1 <=  20'h51986;
               12'b011110111100: data1 <=  20'h61546;
               12'b011110111101: data1 <=  20'h5dd46;
               12'b011110111110: data1 <=  20'h550c9;
               12'b011110111111: data1 <=  20'h520c9;
               12'b011111000000: data1 <=  20'h21908;
               12'b011111000001: data1 <=  20'h70d86;
               12'b011111000010: data1 <=  20'h7a144;
               12'b011111000011: data1 <=  20'h77144;
               12'b011111000100: data1 <=  20'h78643;
               12'b011111000101: data1 <=  20'h5988a;
               12'b011111000110: data1 <=  20'h00306;
               12'b011111000111: data1 <=  20'h064c9;
               12'b011111001000: data1 <=  20'h39686;
               12'b011111001001: data1 <=  20'h5e268;
               12'b011111001010: data1 <=  20'h03946;
               12'b011111001011: data1 <=  20'h3eeae;
               12'b011111001100: data1 <=  20'h41108;
               12'b011111001101: data1 <=  20'h33944;
               12'b011111001110: data1 <=  20'h21c89;
               12'b011111001111: data1 <=  20'h210ca;
               12'b011111010000: data1 <=  20'h1c88d;
               12'b011111010001: data1 <=  20'h1a88d;
               12'b011111010010: data1 <=  20'h2dd26;
               12'b011111010011: data1 <=  20'h26606;
               12'b011111010100: data1 <=  20'h1a60e;
               12'b011111010101: data1 <=  20'h00304;
               12'b011111010110: data1 <=  20'h08926;
               12'b011111010111: data1 <=  20'h075c4;
               12'b011111011000: data1 <=  20'h5a0e9;
               12'b011111011001: data1 <=  20'h14d0a;
               12'b011111011010: data1 <=  20'h14985;
               12'b011111011011: data1 <=  20'h0e88d;
               12'b011111011100: data1 <=  20'h0f473;
               12'b011111011101: data1 <=  20'h2d926;
               12'b011111011110: data1 <=  20'h8aa82;
               12'b011111011111: data1 <=  20'h64304;
               12'b011111100000: data1 <=  20'h14985;
               12'b011111100001: data1 <=  20'h3ed0e;
               12'b011111100010: data1 <=  20'h66cc6;
               12'b011111100011: data1 <=  20'h01958;
               12'b011111100100: data1 <=  20'h211ce;
               12'b011111100101: data1 <=  20'h33d48;
               12'b011111100110: data1 <=  20'h08926;
               12'b011111100111: data1 <=  20'h25b03;
               12'b011111101000: data1 <=  20'h14985;
               12'b011111101001: data1 <=  20'h51ac4;
               12'b011111101010: data1 <=  20'h4d586;
               12'b011111101011: data1 <=  20'h1f526;
               12'b011111101100: data1 <=  20'h1fae6;
               12'b011111101101: data1 <=  20'h25e6c;
               12'b011111101110: data1 <=  20'h088d5;
               12'b011111101111: data1 <=  20'h77a43;
               12'b011111110000: data1 <=  20'h59cc9;
               12'b011111110001: data1 <=  20'h27c8c;
               12'b011111110010: data1 <=  20'h040c9;
               12'b011111110011: data1 <=  20'h008c9;
               12'b011111110100: data1 <=  20'h09896;
               12'b011111110101: data1 <=  20'h3250c;
               12'b011111110110: data1 <=  20'h2f4e9;
               12'b011111110111: data1 <=  20'h4be44;
               12'b011111111000: data1 <=  20'h09896;
               12'b011111111001: data1 <=  20'h08096;
               12'b011111111010: data1 <=  20'h2ce84;
               12'b011111111011: data1 <=  20'h40cc7;
               12'b011111111100: data1 <=  20'h2d944;
               12'b011111111101: data1 <=  20'h12c8f;
               12'b011111111110: data1 <=  20'h03d0c;
               12'b011111111111: data1 <=  20'h0050c;
               12'b100000000000: data1 <=  20'h22cd0;
               12'b100000000001: data1 <=  20'h204d0;
               12'b100000000010: data1 <=  20'h03cd0;
               12'b100000000011: data1 <=  20'h00cd0;
               12'b100000000100: data1 <=  20'h0cb03;
               12'b100000000101: data1 <=  20'h08144;
               12'b100000000110: data1 <=  20'h006e8;
               12'b100000000111: data1 <=  20'h6aa63;
               12'b100000001000: data1 <=  20'h72242;
               12'b100000001001: data1 <=  20'h6a926;
               12'b100000001010: data1 <=  20'h618c9;
               12'b100000001011: data1 <=  20'h5e8c9;
               12'b100000001100: data1 <=  20'h58a86;
               12'b100000001101: data1 <=  20'h3e8ce;
               12'b100000001110: data1 <=  20'h72243;
               12'b100000001111: data1 <=  20'h4c127;
               12'b100000010000: data1 <=  20'h40245;
               12'b100000010001: data1 <=  20'h3ea45;
               12'b100000010010: data1 <=  20'h0d649;
               12'b100000010011: data1 <=  20'h2694a;
               12'b100000010100: data1 <=  20'h5c889;
               12'b100000010101: data1 <=  20'h57889;
               12'b100000010110: data1 <=  20'h09094;
               12'b100000010111: data1 <=  20'h84d83;
               12'b100000011000: data1 <=  20'h09094;
               12'b100000011001: data1 <=  20'h64548;
               12'b100000011010: data1 <=  20'h09094;
               12'b100000011011: data1 <=  20'h00473;
               12'b100000011100: data1 <=  20'h09094;
               12'b100000011101: data1 <=  20'h064c9;
               12'b100000011110: data1 <=  20'h2ca64;
               12'b100000011111: data1 <=  20'h59526;
               12'b100000100000: data1 <=  20'h0a8e6;
               12'b100000100001: data1 <=  20'h015c8;
               12'b100000100010: data1 <=  20'h0a506;
               12'b100000100011: data1 <=  20'h06506;
               12'b100000100100: data1 <=  20'h01a44;
               12'b100000100101: data1 <=  20'h57926;
               12'b100000100110: data1 <=  20'h2ca48;
               12'b100000100111: data1 <=  20'h454c9;
               12'b100000101000: data1 <=  20'h21cc9;
               12'b100000101001: data1 <=  20'h28092;
               12'b100000101010: data1 <=  20'h09094;
               12'b100000101011: data1 <=  20'h08894;
               12'b100000101100: data1 <=  20'h39a46;
               12'b100000101101: data1 <=  20'h1a8c9;
               12'b100000101110: data1 <=  20'h66906;
               12'b100000101111: data1 <=  20'h00248;
               12'b100000110000: data1 <=  20'h20dcc;
               12'b100000110001: data1 <=  20'h13de7;
               12'b100000110010: data1 <=  20'h4e946;
               12'b100000110011: data1 <=  20'h44c8a;
               12'b100000110100: data1 <=  20'h3eec3;
               12'b100000110101: data1 <=  20'h3a4ca;
               12'b100000110110: data1 <=  20'h0fccc;
               12'b100000110111: data1 <=  20'h28092;
               12'b100000111000: data1 <=  20'h33d50;
               12'b100000111001: data1 <=  20'h0850c;
               12'b100000111010: data1 <=  20'h0818e;
               12'b100000111011: data1 <=  20'h58186;
               12'b100000111100: data1 <=  20'h66cc6;
               12'b100000111101: data1 <=  20'h65cc6;
               12'b100000111110: data1 <=  20'h1c48a;
               12'b100000111111: data1 <=  20'h76e63;
               12'b100001000000: data1 <=  20'h350c8;
               12'b100001000001: data1 <=  20'h08516;
               12'b100001000010: data1 <=  20'h350c8;
               12'b100001000011: data1 <=  20'h338c8;
               12'b100001000100: data1 <=  20'h22cc9;
               12'b100001000101: data1 <=  20'h25b04;
               12'b100001000110: data1 <=  20'h4e946;
               12'b100001000111: data1 <=  20'h4b146;
               12'b100001001000: data1 <=  20'h26a63;
               12'b100001001001: data1 <=  20'h25e63;
               12'b100001001010: data1 <=  20'h01209;
               12'b100001001011: data1 <=  20'h06705;
               12'b100001001100: data1 <=  20'h264cf;
               12'b100001001101: data1 <=  20'h27cc9;
               12'b100001001110: data1 <=  20'h6a643;
               12'b100001001111: data1 <=  20'h8b242;
               12'b100001010000: data1 <=  20'h4b8c9;
               12'b100001010001: data1 <=  20'h4f8c9;
               12'b100001010010: data1 <=  20'h4b0c9;
               12'b100001010011: data1 <=  20'h5a48a;
               12'b100001010100: data1 <=  20'h27cd0;
               12'b100001010101: data1 <=  20'h2d94a;
               12'b100001010110: data1 <=  20'h130cd;
               12'b100001010111: data1 <=  20'h0accd;
               12'b100001011000: data1 <=  20'h078c9;
               12'b100001011001: data1 <=  20'h110cb;
               12'b100001011010: data1 <=  20'h0c8cb;
               12'b100001011011: data1 <=  20'h4d5e6;
               12'b100001011100: data1 <=  20'h0d283;
               12'b100001011101: data1 <=  20'h28089;
               12'b100001011110: data1 <=  20'h26d8e;
               12'b100001011111: data1 <=  20'h024c9;
               12'b100001100000: data1 <=  20'h01d26;
               12'b100001100001: data1 <=  20'h280c9;
               12'b100001100010: data1 <=  20'h07594;
               12'b100001100011: data1 <=  20'h2d643;
               12'b100001100100: data1 <=  20'h2be43;
               12'b100001100101: data1 <=  20'h7de43;
               12'b100001100110: data1 <=  20'h27cc9;
               12'b100001100111: data1 <=  20'h0e18f;
               12'b100001101000: data1 <=  20'h13643;
               12'b100001101001: data1 <=  20'h1dc92;
               12'b100001101010: data1 <=  20'h06663;
               12'b100001101011: data1 <=  20'h015e4;
               12'b100001101100: data1 <=  20'h0ddc5;
               12'b100001101101: data1 <=  20'h0cece;
               12'b100001101110: data1 <=  20'h5fcc9;
               12'b100001101111: data1 <=  20'h6be43;
               12'b100001110000: data1 <=  20'h27c72;
               12'b100001110001: data1 <=  20'h00a83;
               12'b100001110010: data1 <=  20'h1a4ac;
               12'b100001110011: data1 <=  20'h27985;
               12'b100001110100: data1 <=  20'h4d4cc;
               12'b100001110101: data1 <=  20'h5b10a;
               12'b100001110110: data1 <=  20'h5810a;
               12'b100001110111: data1 <=  20'h73186;
               12'b100001111000: data1 <=  20'h130c9;
               12'b100001111001: data1 <=  20'h15874;
               12'b100001111010: data1 <=  20'h269c6;
               12'b100001111011: data1 <=  20'h20d8d;
               12'b100001111100: data1 <=  20'h1a48f;
               12'b100001111101: data1 <=  20'h665e4;
               12'b100001111110: data1 <=  20'h33cce;
               12'b100001111111: data1 <=  20'h27546;
               12'b100010000000: data1 <=  20'h1fe43;
               12'b100010000001: data1 <=  20'h079e8;
               12'b100010000010: data1 <=  20'h08112;
               12'b100010000011: data1 <=  20'h3eb03;
               12'b100010000100: data1 <=  20'h0c8cd;
               12'b100010000101: data1 <=  20'h0410a;
               12'b100010000110: data1 <=  20'h07949;
               12'b100010000111: data1 <=  20'h26e43;
               12'b100010001000: data1 <=  20'h06703;
               12'b100010001001: data1 <=  20'h1bccb;
               12'b100010001010: data1 <=  20'h0010a;
               12'b100010001011: data1 <=  20'h65243;
               12'b100010001100: data1 <=  20'h64a43;
               12'b100010001101: data1 <=  20'h00e4a;
               12'b100010001110: data1 <=  20'h13695;
               12'b100010001111: data1 <=  20'h2d5c3;
               12'b100010010000: data1 <=  20'h38586;
               12'b100010010001: data1 <=  20'h586a4;
               12'b100010010010: data1 <=  20'h57aa4;
               12'b100010010011: data1 <=  20'h84a43;
               12'b100010010100: data1 <=  20'h83a43;
               12'b100010010101: data1 <=  20'h1dc92;
               12'b100010010110: data1 <=  20'h2ca43;
               12'b100010010111: data1 <=  20'h1dc92;
               12'b100010011000: data1 <=  20'h5f946;
               12'b100010011001: data1 <=  20'h53969;
               12'b100010011010: data1 <=  20'h2588a;
               12'b100010011011: data1 <=  20'h67d26;
               12'b100010011100: data1 <=  20'h1f892;
               12'b100010011101: data1 <=  20'h3450a;
               12'b100010011110: data1 <=  20'h33d0a;
               12'b100010011111: data1 <=  20'h34585;
               12'b100010100000: data1 <=  20'h33d27;
               12'b100010100001: data1 <=  20'h34585;
               12'b100010100010: data1 <=  20'h27527;
               12'b100010100011: data1 <=  20'h34585;
               12'b100010100100: data1 <=  20'h21c92;
               12'b100010100101: data1 <=  20'h209cc;
               12'b100010100110: data1 <=  20'h06564;
               12'b100010100111: data1 <=  20'h40cca;
               12'b100010101000: data1 <=  20'h6ad66;
               12'b100010101001: data1 <=  20'h67d26;
               12'b100010101010: data1 <=  20'h3ee42;
               12'b100010101011: data1 <=  20'h1a98d;
               12'b100010101100: data1 <=  20'h70a43;
               12'b100010101101: data1 <=  20'h72243;
               12'b100010101110: data1 <=  20'h64126;
               12'b100010101111: data1 <=  20'h61126;
               12'b100010110000: data1 <=  20'h5e526;
               12'b100010110001: data1 <=  20'h098d0;
               12'b100010110010: data1 <=  20'h078d0;
               12'b100010110011: data1 <=  20'h220ca;
               12'b100010110100: data1 <=  20'h210ca;
               12'b100010110101: data1 <=  20'h028d8;
               12'b100010110110: data1 <=  20'h19c94;
               12'b100010110111: data1 <=  20'h038c9;
               12'b100010111000: data1 <=  20'h010c9;
               12'b100010111001: data1 <=  20'h20645;
               12'b100010111010: data1 <=  20'h26cc9;
               12'b100010111011: data1 <=  20'h0e5e8;
               12'b100010111100: data1 <=  20'h0d1e8;
               12'b100010111101: data1 <=  20'h02889;
               12'b100010111110: data1 <=  20'h19ccc;
               12'b100010111111: data1 <=  20'h04112;
               12'b100011000000: data1 <=  20'h00112;
               12'b100011000001: data1 <=  20'h2bf06;
               12'b100011000010: data1 <=  20'h2cdc3;
               12'b100011000011: data1 <=  20'h3490f;
               12'b100011000100: data1 <=  20'h01d4e;
               12'b100011000101: data1 <=  20'h41d0a;
               12'b100011000110: data1 <=  20'h00c89;
               12'b100011000111: data1 <=  20'h0a4c8;
               12'b100011001000: data1 <=  20'h06cc8;
               12'b100011001001: data1 <=  20'h2664c;
               12'b100011001010: data1 <=  20'h4c204;
               12'b100011001011: data1 <=  20'h3960f;
               12'b100011001100: data1 <=  20'h3f50a;
               12'b100011001101: data1 <=  20'h72a06;
               12'b100011001110: data1 <=  20'h64985;
               12'b100011001111: data1 <=  20'h5b124;
               12'b100011010000: data1 <=  20'h59526;
               12'b100011010001: data1 <=  20'h3fa0c;
               12'b100011010010: data1 <=  20'h51666;
               12'b100011010011: data1 <=  20'h53d26;
               12'b100011010100: data1 <=  20'h01477;
               12'b100011010101: data1 <=  20'h32306;
               12'b100011010110: data1 <=  20'h1f4ac;
               12'b100011010111: data1 <=  20'h00e72;
               12'b100011011000: data1 <=  20'h470cc;
               12'b100011011001: data1 <=  20'h1f708;
               12'b100011011010: data1 <=  20'h72124;
               12'b100011011011: data1 <=  20'h34146;
               12'b100011011100: data1 <=  20'h2c683;
               12'b100011011101: data1 <=  20'h030f4;
               12'b100011011110: data1 <=  20'h014f4;
               12'b100011011111: data1 <=  20'h10052;
               12'b100011100000: data1 <=  20'h3354c;
               12'b100011100001: data1 <=  20'h39d88;
               12'b100011100010: data1 <=  20'h2d86e;
               12'b100011100011: data1 <=  20'h0f590;
               12'b100011100100: data1 <=  20'h01cc9;
               12'b100011100101: data1 <=  20'h5ad24;
               12'b100011100110: data1 <=  20'h4b2c4;
               12'b100011100111: data1 <=  20'h4b6c6;
               12'b100011101000: data1 <=  20'h27126;
               12'b100011101001: data1 <=  20'h02889;
               12'b100011101010: data1 <=  20'h32e47;
               12'b100011101011: data1 <=  20'h25b06;
               12'b100011101100: data1 <=  20'h44f0a;
               12'b100011101101: data1 <=  20'h13a55;
               12'b100011101110: data1 <=  20'h4cc8a;
               12'b100011101111: data1 <=  20'h66948;
               12'b100011110000: data1 <=  20'h278c9;
               12'b100011110001: data1 <=  20'h418cc;
               12'b100011110010: data1 <=  20'h400cc;
               12'b100011110011: data1 <=  20'h4f0cc;
               12'b100011110100: data1 <=  20'h4b8cc;
               12'b100011110101: data1 <=  20'h604c9;
               12'b100011110110: data1 <=  20'h5fcc9;
               12'b100011110111: data1 <=  20'h80944;
               12'b100011111000: data1 <=  20'h7d144;
               12'b100011111001: data1 <=  20'h6d126;
               12'b100011111010: data1 <=  20'h0d5c4;
               12'b100011111011: data1 <=  20'h08d44;
               12'b100011111100: data1 <=  20'h5dd44;
               12'b100011111101: data1 <=  20'h11473;
               12'b100011111110: data1 <=  20'h4c128;
               12'b100011111111: data1 <=  20'h2ccac;
               12'b100100000000: data1 <=  20'h06703;
               12'b100100000001: data1 <=  20'h33984;
               12'b100100000010: data1 <=  20'h1788a;
               12'b100100000011: data1 <=  20'h25926;
               12'b100100000100: data1 <=  20'h048d6;
               12'b100100000101: data1 <=  20'h000d6;
               12'b100100000110: data1 <=  20'h5f263;
               12'b100100000111: data1 <=  20'h2e48f;
               12'b100100001000: data1 <=  20'h27cc9;
               12'b100100001001: data1 <=  20'h83643;
               12'b100100001010: data1 <=  20'h1494f;
               12'b100100001011: data1 <=  20'h2c243;
               12'b100100001100: data1 <=  20'h0e926;
               12'b100100001101: data1 <=  20'h3eb0e;
               12'b100100001110: data1 <=  20'h3b90a;
               12'b100100001111: data1 <=  20'h21c89;
               12'b100100010000: data1 <=  20'h3b90a;
               12'b100100010001: data1 <=  20'h4694a;
               12'b100100010010: data1 <=  20'h52644;
               12'b100100010011: data1 <=  20'h00262;
               12'b100100010100: data1 <=  20'h70b06;
               12'b100100010101: data1 <=  20'h1a910;
               12'b100100010110: data1 <=  20'h33d44;
               12'b100100010111: data1 <=  20'h12cc9;
               12'b100100011000: data1 <=  20'h610e9;
               12'b100100011001: data1 <=  20'h71586;
               12'b100100011010: data1 <=  20'h5a8c9;
               12'b100100011011: data1 <=  20'h5e5e8;
               12'b100100011100: data1 <=  20'h27cd0;
               12'b100100011101: data1 <=  20'h270ec;
               12'b100100011110: data1 <=  20'h290c9;
               12'b100100011111: data1 <=  20'h58cc9;
               12'b100100100000: data1 <=  20'h348c9;
               12'b100100100001: data1 <=  20'h27092;
               12'b100100100010: data1 <=  20'h3bccc;
               12'b100100100011: data1 <=  20'h394cc;
               12'b100100100100: data1 <=  20'h61526;
               12'b100100100101: data1 <=  20'h7d244;
               12'b100100100110: data1 <=  20'h73d26;
               12'b100100100111: data1 <=  20'h71126;
               12'b100100101000: data1 <=  20'h65a43;
               12'b100100101001: data1 <=  20'h64243;
               12'b100100101010: data1 <=  20'h11496;
               12'b100100101011: data1 <=  20'h0cc96;
               12'b100100101100: data1 <=  20'h03c58;
               12'b100100101101: data1 <=  20'h7de04;
               12'b100100101110: data1 <=  20'h28492;
               12'b100100101111: data1 <=  20'h3a14e;
               12'b100100110000: data1 <=  20'h290c9;
               12'b100100110001: data1 <=  20'h264e9;
               12'b100100110010: data1 <=  20'h1e094;
               12'b100100110011: data1 <=  20'h274c9;
               12'b100100110100: data1 <=  20'h01d4e;
               12'b100100110101: data1 <=  20'h06e46;
               12'b100100110110: data1 <=  20'h03c58;
               12'b100100110111: data1 <=  20'h01c58;
               12'b100100111000: data1 <=  20'h4e4c7;
               12'b100100111001: data1 <=  20'h4c4c7;
               12'b100100111010: data1 <=  20'h20253;
               12'b100100111011: data1 <=  20'h26d26;
               12'b100100111100: data1 <=  20'h21926;
               12'b100100111101: data1 <=  20'h64d48;
               12'b100100111110: data1 <=  20'h36caf;
               12'b100100111111: data1 <=  20'h320af;
               12'b100101000000: data1 <=  20'h1e094;
               12'b100101000001: data1 <=  20'h19094;
               12'b100101000010: data1 <=  20'h2d944;
               12'b100101000011: data1 <=  20'h77dc4;
               12'b100101000100: data1 <=  20'h47583;
               12'b100101000101: data1 <=  20'h06703;
               12'b100101000110: data1 <=  20'h0e5d4;
               12'b100101000111: data1 <=  20'h514c9;
               12'b100101001000: data1 <=  20'h03493;
               12'b100101001001: data1 <=  20'h451c3;
               12'b100101001010: data1 <=  20'h08214;
               12'b100101001011: data1 <=  20'h3eaa9;
               12'b100101001100: data1 <=  20'h785e5;
               12'b100101001101: data1 <=  20'h408c6;
               12'b100101001110: data1 <=  20'h08214;
               12'b100101001111: data1 <=  20'h06a14;
               12'b100101010000: data1 <=  20'h1d06c;
               12'b100101010001: data1 <=  20'h1a46c;
               12'b100101010010: data1 <=  20'h27548;
               12'b100101010011: data1 <=  20'h394c6;
               12'b100101010100: data1 <=  20'h20d84;
               12'b100101010101: data1 <=  20'h0ecaf;
               12'b100101010110: data1 <=  20'h03d26;
               12'b100101010111: data1 <=  20'h0196a;
               12'b100101011000: data1 <=  20'h2ec8c;
               12'b100101011001: data1 <=  20'h0e524;
               12'b100101011010: data1 <=  20'h019a6;
               12'b100101011011: data1 <=  20'h28092;
               12'b100101011100: data1 <=  20'h348c9;
               12'b100101011101: data1 <=  20'h71546;
               12'b100101011110: data1 <=  20'h58a83;
               12'b100101011111: data1 <=  20'h5e526;
               12'b100101100000: data1 <=  20'h03493;
               12'b100101100001: data1 <=  20'h01c93;
               12'b100101100010: data1 <=  20'h196c2;
               12'b100101100011: data1 <=  20'h00126;
               12'b100101100100: data1 <=  20'h00312;
               12'b100101100101: data1 <=  20'h0d608;
               12'b100101100110: data1 <=  20'h26646;
               12'b100101100111: data1 <=  20'h070ca;
               12'b100101101000: data1 <=  20'h03526;
               12'b100101101001: data1 <=  20'h00926;
               12'b100101101010: data1 <=  20'h0f08f;
               12'b100101101011: data1 <=  20'h018ea;
               12'b100101101100: data1 <=  20'h0d284;
               12'b100101101101: data1 <=  20'h45663;
               12'b100101101110: data1 <=  20'h348c9;
               12'b100101101111: data1 <=  20'h340c9;
               12'b100101110000: data1 <=  20'h35489;
               12'b100101110001: data1 <=  20'h45929;
               12'b100101110010: data1 <=  20'h39245;
               12'b100101110011: data1 <=  20'h19854;
               12'b100101110100: data1 <=  20'h6dd06;
               12'b100101110101: data1 <=  20'h84242;
               12'b100101110110: data1 <=  20'h1a5e6;
               12'b100101110111: data1 <=  20'h5e586;
               12'b100101111000: data1 <=  20'h364c9;
               12'b100101111001: data1 <=  20'h4ba84;
               12'b100101111010: data1 <=  20'h6a706;
               12'b100101111011: data1 <=  20'h65d24;
               12'b100101111100: data1 <=  20'h0a096;
               12'b100101111101: data1 <=  20'h07896;
               12'b100101111110: data1 <=  20'h54109;
               12'b100101111111: data1 <=  20'h07cc9;
               12'b100110000000: data1 <=  20'h1bc72;
               12'b100110000001: data1 <=  20'h33586;
               12'b100110000010: data1 <=  20'h2f8a8;
               12'b100110000011: data1 <=  20'h2cca8;
               12'b100110000100: data1 <=  20'h288cc;
               12'b100110000101: data1 <=  20'h270cc;
               12'b100110000110: data1 <=  20'h399c8;
               12'b100110000111: data1 <=  20'h0886e;
               12'b100110001000: data1 <=  20'h288cc;
               12'b100110001001: data1 <=  20'h20492;
               12'b100110001010: data1 <=  20'h26a12;
               12'b100110001011: data1 <=  20'h1a4f4;
               12'b100110001100: data1 <=  20'h3590c;
               12'b100110001101: data1 <=  20'h40cce;
               12'b100110001110: data1 <=  20'h21926;
               12'b100110001111: data1 <=  20'h1b472;
               12'b100110010000: data1 <=  20'h196ce;
               12'b100110010001: data1 <=  20'h2c642;
               12'b100110010010: data1 <=  20'h288cc;
               12'b100110010011: data1 <=  20'h20d27;
               12'b100110010100: data1 <=  20'h2ec8c;
               12'b100110010101: data1 <=  20'h2dc8c;
               12'b100110010110: data1 <=  20'h0e556;
               12'b100110010111: data1 <=  20'h06474;
               12'b100110011000: data1 <=  20'h52644;
               12'b100110011001: data1 <=  20'h51e44;
               12'b100110011010: data1 <=  20'h61926;
               12'b100110011011: data1 <=  20'h5dd26;
               12'b100110011100: data1 <=  20'h01a58;
               12'b100110011101: data1 <=  20'h270cc;
               12'b100110011110: data1 <=  20'h2dd44;
               12'b100110011111: data1 <=  20'h38a46;
               12'b100110100000: data1 <=  20'h27243;
               12'b100110100001: data1 <=  20'h2d928;
               12'b100110100010: data1 <=  20'h4d8cc;
               12'b100110100011: data1 <=  20'h58643;
               12'b100110100100: data1 <=  20'h6e127;
               12'b100110100101: data1 <=  20'h4b546;
               12'b100110100110: data1 <=  20'h6e127;
               12'b100110100111: data1 <=  20'h15473;
               12'b100110101000: data1 <=  20'h6e127;
               12'b100110101001: data1 <=  20'h07d69;
               12'b100110101010: data1 <=  20'h6e127;
               12'b100110101011: data1 <=  20'h20d66;
               12'b100110101100: data1 <=  20'h2fd05;
               12'b100110101101: data1 <=  20'h19a93;
               12'b100110101110: data1 <=  20'h06ea6;
               12'b100110101111: data1 <=  20'h20d8e;
               12'b100110110000: data1 <=  20'h024c9;
               12'b100110110001: data1 <=  20'h45505;
               12'b100110110010: data1 <=  20'h2fd05;
               12'b100110110011: data1 <=  20'h2bd05;
               12'b100110110100: data1 <=  20'h6e127;
               12'b100110110101: data1 <=  20'h2790a;
               12'b100110110110: data1 <=  20'h61929;
               12'b100110110111: data1 <=  20'h5dd29;
               12'b100110111000: data1 <=  20'h41927;
               12'b100110111001: data1 <=  20'h3f527;
               12'b100110111010: data1 <=  20'h61148;
               12'b100110111011: data1 <=  20'h064cc;
               12'b100110111100: data1 <=  20'h028cc;
               12'b100110111101: data1 <=  20'h01d4c;
               12'b100110111110: data1 <=  20'h07608;
               12'b100110111111: data1 <=  20'h83663;
               12'b100111000000: data1 <=  20'h39e44;
               12'b100111000001: data1 <=  20'h19d26;
               12'b100111000010: data1 <=  20'h088cf;
               12'b100111000011: data1 <=  20'h398c6;
               12'b100111000100: data1 <=  20'h079c9;
               12'b100111000101: data1 <=  20'h00d14;
               12'b100111000110: data1 <=  20'h014e9;
               12'b100111000111: data1 <=  20'h27185;
               12'b100111001000: data1 <=  20'h0650e;
               12'b100111001001: data1 <=  20'h4bac4;
               12'b100111001010: data1 <=  20'h6c4c6;
               12'b100111001011: data1 <=  20'h0acc7;
               12'b100111001100: data1 <=  20'h000c6;
               12'b100111001101: data1 <=  20'h26a32;
               12'b100111001110: data1 <=  20'h01986;
               12'b100111001111: data1 <=  20'h2ce44;
               12'b100111010000: data1 <=  20'h4c146;
               12'b100111010001: data1 <=  20'h3a14c;
               12'b100111010010: data1 <=  20'h06703;
               12'b100111010011: data1 <=  20'h480c6;
               12'b100111010100: data1 <=  20'h460c6;
               12'b100111010101: data1 <=  20'h3f663;
               12'b100111010110: data1 <=  20'h0c8c9;
               12'b100111010111: data1 <=  20'h67946;
               12'b100111011000: data1 <=  20'h64146;
               12'b100111011001: data1 <=  20'h54d26;
               12'b100111011010: data1 <=  20'h64243;
               12'b100111011011: data1 <=  20'h65a43;
               12'b100111011100: data1 <=  20'h70926;
               12'b100111011101: data1 <=  20'h54d26;
               12'b100111011110: data1 <=  20'h0e0c9;
               12'b100111011111: data1 <=  20'h35c8c;
               12'b100111100000: data1 <=  20'h53508;
               12'b100111100001: data1 <=  20'h7e243;
               12'b100111100010: data1 <=  20'h3348c;
               12'b100111100011: data1 <=  20'h2d983;
               12'b100111100100: data1 <=  20'h28089;
               12'b100111100101: data1 <=  20'h7e643;
               12'b100111100110: data1 <=  20'h7d643;
               12'b100111100111: data1 <=  20'h0acd4;
               12'b100111101000: data1 <=  20'h064d4;
               12'b100111101001: data1 <=  20'h16092;
               12'b100111101010: data1 <=  20'h0c8cc;
               12'b100111101011: data1 <=  20'h3b586;
               12'b100111101100: data1 <=  20'h14892;
               12'b100111101101: data1 <=  20'h038c9;
               12'b100111101110: data1 <=  20'h38586;
               12'b100111101111: data1 <=  20'h1c914;
               12'b100111110000: data1 <=  20'h19914;
               12'b100111110001: data1 <=  20'h54d26;
               12'b100111110010: data1 <=  20'h51926;
               12'b100111110011: data1 <=  20'h5ea43;
               12'b100111110100: data1 <=  20'h52926;
               12'b100111110101: data1 <=  20'h01643;
               12'b100111110110: data1 <=  20'h0e8c7;
               12'b100111110111: data1 <=  20'h08926;
               12'b100111111000: data1 <=  20'h07d26;
               12'b100111111001: data1 <=  20'h26dc6;
               12'b100111111010: data1 <=  20'h0e8cd;
               12'b100111111011: data1 <=  20'h46586;
               12'b100111111100: data1 <=  20'h0724f;
               12'b100111111101: data1 <=  20'h034c7;
               12'b100111111110: data1 <=  20'h13a06;
               12'b100111111111: data1 <=  20'h0946c;
               12'b101000000000: data1 <=  20'h2d8c9;
               12'b101000000001: data1 <=  20'h03498;
               12'b101000000010: data1 <=  20'h01c98;
               12'b101000000011: data1 <=  20'h3b0ac;
               12'b101000000100: data1 <=  20'h5f926;
               12'b101000000101: data1 <=  20'h2d246;
               12'b101000000110: data1 <=  20'h3a4ac;
               12'b101000000111: data1 <=  20'h6b626;
               12'b101000001000: data1 <=  20'h12e4e;
               12'b101000001001: data1 <=  20'h06702;
               12'b101000001010: data1 <=  20'h5de43;
               12'b101000001011: data1 <=  20'h024c9;
               12'b101000001100: data1 <=  20'h139cc;
               12'b101000001101: data1 <=  20'h0946c;
               12'b101000001110: data1 <=  20'h020c9;
               12'b101000001111: data1 <=  20'h280ca;
               12'b101000010000: data1 <=  20'h014c9;
               12'b101000010001: data1 <=  20'h00aa7;
               12'b101000010010: data1 <=  20'h46585;
               12'b101000010011: data1 <=  20'h2dd28;
               12'b101000010100: data1 <=  20'h27cd2;
               12'b101000010101: data1 <=  20'h5b50a;
               12'b101000010110: data1 <=  20'h57d0a;
               12'b101000010111: data1 <=  20'h02d0a;
               12'b101000011000: data1 <=  20'h0150a;
               12'b101000011001: data1 <=  20'h07d85;
               12'b101000011010: data1 <=  20'h4b642;
               12'b101000011011: data1 <=  20'h32a86;
               12'b101000011100: data1 <=  20'h27527;
               12'b101000011101: data1 <=  20'h21d10;
               12'b101000011110: data1 <=  20'h39208;
               12'b101000011111: data1 <=  20'h33d44;
               12'b101000100000: data1 <=  20'h4cd48;
               12'b101000100001: data1 <=  20'h791e4;
               12'b101000100010: data1 <=  20'h00649;
               12'b101000100011: data1 <=  20'h1c548;
               12'b101000100100: data1 <=  20'h64e44;
               12'b101000100101: data1 <=  20'h2dd4c;
               12'b101000100110: data1 <=  20'h2d54c;
               12'b101000100111: data1 <=  20'h26a47;
               12'b101000101000: data1 <=  20'h6a643;
               12'b101000101001: data1 <=  20'h6b243;
               12'b101000101010: data1 <=  20'h198ca;
               12'b101000101011: data1 <=  20'h04118;
               12'b101000101100: data1 <=  20'h0110f;
               12'b101000101101: data1 <=  20'h04118;
               12'b101000101110: data1 <=  20'h19649;
               12'b101000101111: data1 <=  20'h4ed26;
               12'b101000110000: data1 <=  20'h39246;
               12'b101000110001: data1 <=  20'h23cc9;
               12'b101000110010: data1 <=  20'h1f4c9;
               12'b101000110011: data1 <=  20'h2ce44;
               12'b101000110100: data1 <=  20'h06d94;
               12'b101000110101: data1 <=  20'h044d7;
               12'b101000110110: data1 <=  20'h25c52;
               12'b101000110111: data1 <=  20'h34146;
               12'b101000111000: data1 <=  20'h25a86;
               12'b101000111001: data1 <=  20'h4dd85;
               12'b101000111010: data1 <=  20'h19073;
               12'b101000111011: data1 <=  20'h0b072;
               12'b101000111100: data1 <=  20'h06c72;
               12'b101000111101: data1 <=  20'h3f643;
               12'b101000111110: data1 <=  20'h1a149;
               12'b101000111111: data1 <=  20'h531c7;
               12'b101001000000: data1 <=  20'h521c7;
               12'b101001000001: data1 <=  20'h5fd26;
               12'b101001000010: data1 <=  20'h5890a;
               12'b101001000011: data1 <=  20'h5a08a;
               12'b101001000100: data1 <=  20'h32cb0;
               12'b101001000101: data1 <=  20'h42526;
               12'b101001000110: data1 <=  20'h3e926;
               12'b101001000111: data1 <=  20'h2d589;
               12'b101001001000: data1 <=  20'h40ca8;
               12'b101001001001: data1 <=  20'h0946c;
               12'b101001001010: data1 <=  20'h5fcc9;
               12'b101001001011: data1 <=  20'h298e6;
               12'b101001001100: data1 <=  20'h08496;
               12'b101001001101: data1 <=  20'h271c3;
               12'b101001001110: data1 <=  20'h70a63;
               12'b101001001111: data1 <=  20'h044d8;
               12'b101001010000: data1 <=  20'h515e6;
               12'b101001010001: data1 <=  20'h27d4e;
               12'b101001010010: data1 <=  20'h25d0a;
               12'b101001010011: data1 <=  20'h27585;
               12'b101001010100: data1 <=  20'h2d926;
               12'b101001010101: data1 <=  20'h33dce;
               12'b101001010110: data1 <=  20'h32dce;
               12'b101001010111: data1 <=  20'h345a4;
               12'b101001011000: data1 <=  20'h0d4cc;
               12'b101001011001: data1 <=  20'h40226;
               12'b101001011010: data1 <=  20'h3ee26;
               12'b101001011011: data1 <=  20'h2fd09;
               12'b101001011100: data1 <=  20'h2bd09;
               12'b101001011101: data1 <=  20'h3870a;
               12'b101001011110: data1 <=  20'h0d5e8;
               12'b101001011111: data1 <=  20'h0da48;
               12'b101001100000: data1 <=  20'h06644;
               12'b101001100001: data1 <=  20'h11872;
               12'b101001100010: data1 <=  20'h13073;
               12'b101001100011: data1 <=  20'h368d0;
               12'b101001100100: data1 <=  20'h320d0;
               12'b101001100101: data1 <=  20'h72966;
               12'b101001100110: data1 <=  20'h26985;
               12'b101001100111: data1 <=  20'h27585;
               12'b101001101000: data1 <=  20'h14526;
               12'b101001101001: data1 <=  20'h27585;
               12'b101001101010: data1 <=  20'h344c7;
               12'b101001101011: data1 <=  20'h0e926;
               12'b101001101100: data1 <=  20'h598c9;
               12'b101001101101: data1 <=  20'h0e926;
               12'b101001101110: data1 <=  20'h13e14;
               12'b101001101111: data1 <=  20'h2754c;
               12'b101001110000: data1 <=  20'h0c8ec;
               12'b101001110001: data1 <=  20'h6d566;
               12'b101001110010: data1 <=  20'h2cd88;
               12'b101001110011: data1 <=  20'h46d0a;
               12'b101001110100: data1 <=  20'h08889;
               12'b101001110101: data1 <=  20'h03876;
               12'b101001110110: data1 <=  20'h01c76;
               12'b101001110111: data1 <=  20'h2ce44;
               12'b101001111000: data1 <=  20'h0f08f;
               12'b101001111001: data1 <=  20'h0946c;
               12'b101001111010: data1 <=  20'h0024d;
               12'b101001111011: data1 <=  20'h04078;
               12'b101001111100: data1 <=  20'h01478;
               12'b101001111101: data1 <=  20'h604a8;
               12'b101001111110: data1 <=  20'h71242;
               12'b101001111111: data1 <=  20'h32a83;
               12'b101010000000: data1 <=  20'h27526;
               12'b101010000001: data1 <=  20'h0d66a;
               12'b101010000010: data1 <=  20'h2c663;
               12'b101010000011: data1 <=  20'h29524;
               12'b101010000100: data1 <=  20'h0d248;
               12'b101010000101: data1 <=  20'h3adc4;
               12'b101010000110: data1 <=  20'h1a0d0;
               12'b101010000111: data1 <=  20'h35d30;
               12'b101010001000: data1 <=  20'h32130;
               12'b101010001001: data1 <=  20'h048ce;
               12'b101010001010: data1 <=  20'h000ce;
               12'b101010001011: data1 <=  20'h03cd6;
               12'b101010001100: data1 <=  20'h00cd6;
               12'b101010001101: data1 <=  20'h0f994;
               12'b101010001110: data1 <=  20'h0c994;
               12'b101010001111: data1 <=  20'h28489;
               12'b101010010000: data1 <=  20'h024d0;
               12'b101010010001: data1 <=  20'h0946c;
               12'b101010010010: data1 <=  20'h19e46;
               12'b101010010011: data1 <=  20'h20a08;
               12'b101010010100: data1 <=  20'h51546;
               12'b101010010101: data1 <=  20'h59926;
               12'b101010010110: data1 <=  20'h0e126;
               12'b101010010111: data1 <=  20'h09d48;
               12'b101010011000: data1 <=  20'h0886c;
               12'b101010011001: data1 <=  20'h1a989;
               12'b101010011010: data1 <=  20'h20d86;
               12'b101010011011: data1 <=  20'h06905;
               12'b101010011100: data1 <=  20'h4e0c8;
               12'b101010011101: data1 <=  20'h4bd86;
               12'b101010011110: data1 <=  20'h72d86;
               12'b101010011111: data1 <=  20'h524c6;
               12'b101010100000: data1 <=  20'h158f2;
               12'b101010100001: data1 <=  20'h39243;
               12'b101010100010: data1 <=  20'h14262;
               12'b101010100011: data1 <=  20'h0d986;
               12'b101010100100: data1 <=  20'h27cc9;
               12'b101010100101: data1 <=  20'h278c9;
               12'b101010100110: data1 <=  20'h3c4af;
               12'b101010100111: data1 <=  20'h390af;
               12'b101010101000: data1 <=  20'h271c6;
               12'b101010101001: data1 <=  20'h2786e;
               12'b101010101010: data1 <=  20'h64305;
               12'b101010101011: data1 <=  20'h7d283;
               12'b101010101100: data1 <=  20'h3fe42;
               12'b101010101101: data1 <=  20'h258ca;
               12'b101010101110: data1 <=  20'h06e83;
               12'b101010101111: data1 <=  20'h538cb;
               12'b101010110000: data1 <=  20'h600c8;
               12'b101010110001: data1 <=  20'h4d4c9;
               12'b101010110010: data1 <=  20'h46242;
               12'b101010110011: data1 <=  20'h261e6;
               12'b101010110100: data1 <=  20'h01a43;
               12'b101010110101: data1 <=  20'h01472;
               12'b101010110110: data1 <=  20'h174ca;
               12'b101010110111: data1 <=  20'h12cca;
               12'b101010111000: data1 <=  20'h21d09;
               12'b101010111001: data1 <=  20'h20d09;
               12'b101010111010: data1 <=  20'h0d683;
               12'b101010111011: data1 <=  20'h0dda4;
               12'b101010111100: data1 <=  20'h044ee;
               12'b101010111101: data1 <=  20'h000ee;
               12'b101010111110: data1 <=  20'h47146;
               12'b101010111111: data1 <=  20'h46146;
               12'b101011000000: data1 <=  20'h28472;
               12'b101011000001: data1 <=  20'h64243;
               12'b101011000010: data1 <=  20'h65a43;
               12'b101011000011: data1 <=  20'h2692a;
               12'b101011000100: data1 <=  20'h2e1e4;
               12'b101011000101: data1 <=  20'h26d86;
               12'b101011000110: data1 <=  20'h07d89;
               12'b101011000111: data1 <=  20'h3a0cc;
               12'b101011001000: data1 <=  20'h221a6;
               12'b101011001001: data1 <=  20'h452cd;
               12'b101011001010: data1 <=  20'h368c6;
               12'b101011001011: data1 <=  20'h320c6;
               12'b101011001100: data1 <=  20'h25b03;
               12'b101011001101: data1 <=  20'h1f546;
               12'b101011001110: data1 <=  20'h2d643;
               12'b101011001111: data1 <=  20'h00146;
               12'b101011010000: data1 <=  20'h04c73;
               12'b101011010001: data1 <=  20'h26990;
               12'b101011010010: data1 <=  20'h2a492;
               12'b101011010011: data1 <=  20'h25c92;
               12'b101011010100: data1 <=  20'h84243;
               12'b101011010101: data1 <=  20'h76d24;
               12'b101011010110: data1 <=  20'h73986;
               12'b101011010111: data1 <=  20'h72524;
               12'b101011011000: data1 <=  20'h67148;
               12'b101011011001: data1 <=  20'h64948;
               12'b101011011010: data1 <=  20'h0394c;
               12'b101011011011: data1 <=  20'h0014c;
               12'b101011011100: data1 <=  20'h5b526;
               12'b101011011101: data1 <=  20'h57926;
               12'b101011011110: data1 <=  20'h5b146;
               12'b101011011111: data1 <=  20'h57946;
               12'b101011100000: data1 <=  20'h71e42;
               12'b101011100001: data1 <=  20'h70a43;
               12'b101011100010: data1 <=  20'h2024c;
               12'b101011100011: data1 <=  20'h140e9;
               12'b101011100100: data1 <=  20'h0126f;
               12'b101011100101: data1 <=  20'h00e04;
               12'b101011100110: data1 <=  20'h4c20c;
               12'b101011100111: data1 <=  20'h13d8f;
               12'b101011101000: data1 <=  20'h1d053;
               12'b101011101001: data1 <=  20'h1a853;
               12'b101011101010: data1 <=  20'h5ad0a;
               12'b101011101011: data1 <=  20'h5850a;
               12'b101011101100: data1 <=  20'h28872;
               12'b101011101101: data1 <=  20'h46186;
               12'b101011101110: data1 <=  20'h21d0a;
               12'b101011101111: data1 <=  20'h1a98a;
               12'b101011110000: data1 <=  20'h33a4a;
               12'b101011110001: data1 <=  20'h3224a;
               12'b101011110010: data1 <=  20'h28872;
               12'b101011110011: data1 <=  20'h57a43;
               12'b101011110100: data1 <=  20'h28872;
               12'b101011110101: data1 <=  20'h27c72;
               12'b101011110110: data1 <=  20'h59243;
               12'b101011110111: data1 <=  20'h1f643;
               12'b101011111000: data1 <=  20'h1fec3;
               12'b101011111001: data1 <=  20'h002aa;
               12'b101011111010: data1 <=  20'h14651;
               12'b101011111011: data1 <=  20'h12e51;
               12'b101011111100: data1 <=  20'h4b30b;
               12'b101011111101: data1 <=  20'h3fa06;
               12'b101011111110: data1 <=  20'h350c8;
               12'b101011111111: data1 <=  20'h59107;
               12'b101100000000: data1 <=  20'h424ce;
               12'b101100000001: data1 <=  20'h3f4ce;
               12'b101100000010: data1 <=  20'h4ca42;
               12'b101100000011: data1 <=  20'h33546;
               12'b101100000100: data1 <=  20'h47d24;
               12'b101100000101: data1 <=  20'h44d26;
               12'b101100000110: data1 <=  20'h0f472;
               12'b101100000111: data1 <=  20'h0f072;
               12'b101100001000: data1 <=  20'h4d4ca;
               12'b101100001001: data1 <=  20'h3ecc9;
               12'b101100001010: data1 <=  20'h39e06;
               12'b101100001011: data1 <=  20'h32526;
               12'b101100001100: data1 <=  20'h2da06;
               12'b101100001101: data1 <=  20'h00243;
               12'b101100001110: data1 <=  20'h028c9;
               12'b101100001111: data1 <=  20'h218c6;
               12'b101100010000: data1 <=  20'h28092;
               12'b101100010001: data1 <=  20'h020c9;
               12'b101100010010: data1 <=  20'h088c9;
               12'b101100010011: data1 <=  20'h00649;
               12'b101100010100: data1 <=  20'h12f03;
               12'b101100010101: data1 <=  20'h59124;
               12'b101100010110: data1 <=  20'h3a50a;
               12'b101100010111: data1 <=  20'h0dda9;
               12'b101100011000: data1 <=  20'h1a209;
               12'b101100011001: data1 <=  20'h1a1c9;
               12'b101100011010: data1 <=  20'h21526;
               12'b101100011011: data1 <=  20'h2c206;
               12'b101100011100: data1 <=  20'h21da9;
               12'b101100011101: data1 <=  20'h1f9a9;
               12'b101100011110: data1 <=  20'h19306;
               12'b101100011111: data1 <=  20'h57d49;
               12'b101100100000: data1 <=  20'h6ba43;
               12'b101100100001: data1 <=  20'h64243;
               12'b101100100010: data1 <=  20'h6c926;
               12'b101100100011: data1 <=  20'h7d6c4;
               12'b101100100100: data1 <=  20'h59906;
               12'b101100100101: data1 <=  20'h2790f;
               12'b101100100110: data1 <=  20'h1a643;
               12'b101100100111: data1 <=  20'h150aa;
               12'b101100101000: data1 <=  20'h33983;
               12'b101100101001: data1 <=  20'h26246;
               12'b101100101010: data1 <=  20'h28092;
               12'b101100101011: data1 <=  20'h210c6;
               12'b101100101100: data1 <=  20'h22c52;
               12'b101100101101: data1 <=  20'h21452;
               12'b101100101110: data1 <=  20'h0ed46;
               12'b101100101111: data1 <=  20'h0724c;
               12'b101100110000: data1 <=  20'h0de36;
               12'b101100110001: data1 <=  20'h01186;
               12'b101100110010: data1 <=  20'h39e06;
               12'b101100110011: data1 <=  20'h024b2;
               12'b101100110100: data1 <=  20'h030c9;
               12'b101100110101: data1 <=  20'h018c9;
               12'b101100110110: data1 <=  20'h088cc;
               12'b101100110111: data1 <=  20'h399a4;
               12'b101100111000: data1 <=  20'h33663;
               12'b101100111001: data1 <=  20'h3a8c8;
               12'b101100111010: data1 <=  20'h3b08f;
               12'b101100111011: data1 <=  20'h008ce;
               12'b101100111100: data1 <=  20'h0a0ce;
               12'b101100111101: data1 <=  20'h070ce;
               12'b101100111110: data1 <=  20'h7de44;
               12'b101100111111: data1 <=  20'h01494;
               12'b101101000000: data1 <=  20'h3610c;
               12'b101101000001: data1 <=  20'h3210c;
               12'b101101000010: data1 <=  20'h54948;
               12'b101101000011: data1 <=  20'h51948;
               12'b101101000100: data1 <=  20'h35c8f;
               12'b101101000101: data1 <=  20'h3348f;
               12'b101101000110: data1 <=  20'h4660c;
               12'b101101000111: data1 <=  20'h4560c;
               12'b101101001000: data1 <=  20'h4e8e9;
               12'b101101001001: data1 <=  20'h08c75;
               12'b101101001010: data1 <=  20'h48124;
               12'b101101001011: data1 <=  20'h3f629;
               12'b101101001100: data1 <=  20'h3550f;
               12'b101101001101: data1 <=  20'h32d0f;
               12'b101101001110: data1 <=  20'h5a548;
               12'b101101001111: data1 <=  20'h70ac6;
               12'b101101010000: data1 <=  20'h64304;
               12'b101101010001: data1 <=  20'h7e983;
               12'b101101010010: data1 <=  20'h4f8cc;
               12'b101101010011: data1 <=  20'h4b0cc;
               12'b101101010100: data1 <=  20'h6e126;
               12'b101101010101: data1 <=  20'h25eca;
               12'b101101010110: data1 <=  20'h6e126;
               12'b101101010111: data1 <=  20'h70a42;
               12'b101101011000: data1 <=  20'h5ea63;
               12'b101101011001: data1 <=  20'h51643;
               12'b101101011010: data1 <=  20'h6e126;
               12'b101101011011: data1 <=  20'h6a526;
               12'b101101011100: data1 <=  20'h6d526;
               12'b101101011101: data1 <=  20'h6b126;
               12'b101101011110: data1 <=  20'h10874;
               12'b101101011111: data1 <=  20'h51708;
               12'b101101100000: data1 <=  20'h088d6;
               default: data1 <= 0;
           endcase
        end

endmodule: rect0_rom
