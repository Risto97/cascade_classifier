module rect1_rom
  #(
     W_DATA = 20,
     DEPTH = 2913,
     W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input ena,
     input [W_ADDR-1:0] addra,
     output [W_DATA-1:0] doa
    );

     logic [W_DATA-1:0] mem [DEPTH-1:0];

     always_ff @(posedge clk)
        begin
           if(ena)
              doa = mem[addra];
        end

     initial begin
         mem[0] =  20'h2d583;
         mem[1] =  20'h1b887;
         mem[2] =  20'h4be43;
         mem[3] =  20'h7f122;
         mem[4] =  20'h20853;
         mem[5] =  20'h52d88;
         mem[6] =  20'h46183;
         mem[7] =  20'h79885;
         mem[8] =  20'h13ce3;
         mem[9] =  20'h33982;
         mem[10] =  20'h1b887;
         mem[11] =  20'h4b664;
         mem[12] =  20'h0e903;
         mem[13] =  20'h59cc5;
         mem[14] =  20'h461c5;
         mem[15] =  20'h141c3;
         mem[16] =  20'h48c66;
         mem[17] =  20'h2184a;
         mem[18] =  20'h3504a;
         mem[19] =  20'h20449;
         mem[20] =  20'h0504b;
         mem[21] =  20'h2790d;
         mem[22] =  20'h28449;
         mem[23] =  20'h7ed42;
         mem[24] =  20'h529c6;
         mem[25] =  20'h14d03;
         mem[26] =  20'h461e3;
         mem[27] =  20'h538a7;
         mem[28] =  20'h2204a;
         mem[29] =  20'h4c866;
         mem[30] =  20'h858c3;
         mem[31] =  20'h335a2;
         mem[32] =  20'h0ac6f;
         mem[33] =  20'h0746f;
         mem[34] =  20'h3410f;
         mem[35] =  20'h26ce6;
         mem[36] =  20'h64aa4;
         mem[37] =  20'h08c4a;
         mem[38] =  20'h51d4a;
         mem[39] =  20'h06c4d;
         mem[40] =  20'h1184d;
         mem[41] =  20'h22173;
         mem[42] =  20'h1e049;
         mem[43] =  20'h1344b;
         mem[44] =  20'h09449;
         mem[45] =  20'h2be61;
         mem[46] =  20'h09449;
         mem[47] =  20'h08c49;
         mem[48] =  20'h224e7;
         mem[49] =  20'h45241;
         mem[50] =  20'h5584b;
         mem[51] =  20'h2bcc3;
         mem[52] =  20'h2d583;
         mem[53] =  20'h21c86;
         mem[54] =  20'h08505;
         mem[55] =  20'h4c242;
         mem[56] =  20'h6acc3;
         mem[57] =  20'h1784d;
         mem[58] =  20'h1384d;
         mem[59] =  20'h08517;
         mem[60] =  20'h45104;
         mem[61] =  20'h5b067;
         mem[62] =  20'h4bd03;
         mem[63] =  20'h33982;
         mem[64] =  20'h534c6;
         mem[65] =  20'h6e122;
         mem[66] =  20'h70e41;
         mem[67] =  20'h3fa06;
         mem[68] =  20'h06c54;
         mem[69] =  20'h07241;
         mem[70] =  20'h1f947;
         mem[71] =  20'h4c5c4;
         mem[72] =  20'h6b0e3;
         mem[73] =  20'h6dd22;
         mem[74] =  20'h6a922;
         mem[75] =  20'h29485;
         mem[76] =  20'h208e7;
         mem[77] =  20'h02885;
         mem[78] =  20'h150c3;
         mem[79] =  20'h28449;
         mem[80] =  20'h02449;
         mem[81] =  20'h28849;
         mem[82] =  20'h28049;
         mem[83] =  20'h344c4;
         mem[84] =  20'h14583;
         mem[85] =  20'h02106;
         mem[86] =  20'h45e04;
         mem[87] =  20'h28466;
         mem[88] =  20'h7f103;
         mem[89] =  20'h28449;
         mem[90] =  20'h538a4;
         mem[91] =  20'h28449;
         mem[92] =  20'h28449;
         mem[93] =  20'h72cc6;
         mem[94] =  20'h90241;
         mem[95] =  20'h4d885;
         mem[96] =  20'h4c905;
         mem[97] =  20'h33d42;
         mem[98] =  20'h64142;
         mem[99] =  20'h78641;
         mem[100] =  20'h0cec1;
         mem[101] =  20'h6be41;
         mem[102] =  20'h1a46f;
         mem[103] =  20'h1e04a;
         mem[104] =  20'h1984a;
         mem[105] =  20'h67143;
         mem[106] =  20'h4c089;
         mem[107] =  20'h03849;
         mem[108] =  20'h40866;
         mem[109] =  20'h364c3;
         mem[110] =  20'h320c3;
         mem[111] =  20'h03849;
         mem[112] =  20'h02049;
         mem[113] =  20'h66122;
         mem[114] =  20'h70922;
         mem[115] =  20'h3504a;
         mem[116] =  20'h790c3;
         mem[117] =  20'h45681;
         mem[118] =  20'h38d26;
         mem[119] =  20'h00d38;
         mem[120] =  20'h26ce5;
         mem[121] =  20'h22ca6;
         mem[122] =  20'h204c6;
         mem[123] =  20'h5ee41;
         mem[124] =  20'h6bd04;
         mem[125] =  20'h77a43;
         mem[126] =  20'h00c66;
         mem[127] =  20'h28092;
         mem[128] =  20'h0844e;
         mem[129] =  20'h13a61;
         mem[130] =  20'h3516d;
         mem[131] =  20'h46d62;
         mem[132] =  20'h4c4aa;
         mem[133] =  20'h68086;
         mem[134] =  20'h65086;
         mem[135] =  20'h240a4;
         mem[136] =  20'h0e904;
         mem[137] =  20'h40182;
         mem[138] =  20'h21c66;
         mem[139] =  20'h7f4c3;
         mem[140] =  20'h4b2c5;
         mem[141] =  20'h1a223;
         mem[142] =  20'h2184a;
         mem[143] =  20'h0ac68;
         mem[144] =  20'h07067;
         mem[145] =  20'h04876;
         mem[146] =  20'h00c76;
         mem[147] =  20'h2fc90;
         mem[148] =  20'h4ba62;
         mem[149] =  20'h538c4;
         mem[150] =  20'h6ae22;
         mem[151] =  20'h5b067;
         mem[152] =  20'h26c85;
         mem[153] =  20'h3686b;
         mem[154] =  20'h32c6b;
         mem[155] =  20'h5fd49;
         mem[156] =  20'h59467;
         mem[157] =  20'h59908;
         mem[158] =  20'h4112e;
         mem[159] =  20'h614c3;
         mem[160] =  20'h01ca8;
         mem[161] =  20'h03466;
         mem[162] =  20'h15d04;
         mem[163] =  20'h03466;
         mem[164] =  20'h06942;
         mem[165] =  20'h03466;
         mem[166] =  20'h02066;
         mem[167] =  20'h7f142;
         mem[168] =  20'h14c49;
         mem[169] =  20'h21182;
         mem[170] =  20'h44e41;
         mem[171] =  20'h452c1;
         mem[172] =  20'h47088;
         mem[173] =  20'h47c66;
         mem[174] =  20'h47066;
         mem[175] =  20'h4cd62;
         mem[176] =  20'h51582;
         mem[177] =  20'h1c566;
         mem[178] =  20'h03151;
         mem[179] =  20'h03838;
         mem[180] =  20'h02438;
         mem[181] =  20'h09c36;
         mem[182] =  20'h08836;
         mem[183] =  20'h2a032;
         mem[184] =  20'h65922;
         mem[185] =  20'h67522;
         mem[186] =  20'h77a41;
         mem[187] =  20'h1c489;
         mem[188] =  20'h70a41;
         mem[189] =  20'h0e0c4;
         mem[190] =  20'h465c3;
         mem[191] =  20'h21c66;
         mem[192] =  20'h53cc8;
         mem[193] =  20'h1a070;
         mem[194] =  20'h14243;
         mem[195] =  20'h790a4;
         mem[196] =  20'h05049;
         mem[197] =  20'h06e41;
         mem[198] =  20'h91261;
         mem[199] =  20'h00849;
         mem[200] =  20'h4c666;
         mem[201] =  20'h06c49;
         mem[202] =  20'h228e6;
         mem[203] =  20'h0ca81;
         mem[204] =  20'h132c1;
         mem[205] =  20'h454e3;
         mem[206] =  20'h4e562;
         mem[207] =  20'h4b162;
         mem[208] =  20'h2e84b;
         mem[209] =  20'h08c66;
         mem[210] =  20'h2e885;
         mem[211] =  20'h40186;
         mem[212] =  20'h2a0c5;
         mem[213] =  20'h64e41;
         mem[214] =  20'h368c3;
         mem[215] =  20'h1f903;
         mem[216] =  20'h03449;
         mem[217] =  20'h19187;
         mem[218] =  20'h0344d;
         mem[219] =  20'h0244d;
         mem[220] =  20'h28c49;
         mem[221] =  20'h2e449;
         mem[222] =  20'h7a122;
         mem[223] =  20'h710e3;
         mem[224] =  20'h73922;
         mem[225] =  20'h7e4a4;
         mem[226] =  20'h614a9;
         mem[227] =  20'h26a02;
         mem[228] =  20'h33d42;
         mem[229] =  20'h58caa;
         mem[230] =  20'h3b4a7;
         mem[231] =  20'h27c49;
         mem[232] =  20'h2ca41;
         mem[233] =  20'h44e41;
         mem[234] =  20'h67122;
         mem[235] =  20'h268e3;
         mem[236] =  20'h03432;
         mem[237] =  20'h02832;
         mem[238] =  20'h2e4aa;
         mem[239] =  20'h7f0e4;
         mem[240] =  20'h5a0a9;
         mem[241] =  20'h0c983;
         mem[242] =  20'h09564;
         mem[243] =  20'h13de3;
         mem[244] =  20'h02113;
         mem[245] =  20'h86123;
         mem[246] =  20'h2e0a4;
         mem[247] =  20'h2e4a4;
         mem[248] =  20'h37068;
         mem[249] =  20'h5e142;
         mem[250] =  20'h6dd42;
         mem[251] =  20'h13a03;
         mem[252] =  20'h488e5;
         mem[253] =  20'h0904d;
         mem[254] =  20'h10c6e;
         mem[255] =  20'h584c5;
         mem[256] =  20'h33d42;
         mem[257] =  20'h0d86e;
         mem[258] =  20'h348a4;
         mem[259] =  20'h6c505;
         mem[260] =  20'h488a4;
         mem[261] =  20'h07066;
         mem[262] =  20'h670c3;
         mem[263] =  20'h658c3;
         mem[264] =  20'h5b068;
         mem[265] =  20'h57da2;
         mem[266] =  20'h09849;
         mem[267] =  20'h02866;
         mem[268] =  20'h0f869;
         mem[269] =  20'h0ec69;
         mem[270] =  20'h7e982;
         mem[271] =  20'h27c49;
         mem[272] =  20'h2d8c3;
         mem[273] =  20'h40907;
         mem[274] =  20'h33d44;
         mem[275] =  20'h190c3;
         mem[276] =  20'h10434;
         mem[277] =  20'h258c3;
         mem[278] =  20'h16835;
         mem[279] =  20'h02037;
         mem[280] =  20'h42522;
         mem[281] =  20'h3e922;
         mem[282] =  20'h66122;
         mem[283] =  20'h64122;
         mem[284] =  20'h40cc4;
         mem[285] =  20'h02113;
         mem[286] =  20'h2e106;
         mem[287] =  20'h2884a;
         mem[288] =  20'h3b4a6;
         mem[289] =  20'h01833;
         mem[290] =  20'h0404a;
         mem[291] =  20'h00866;
         mem[292] =  20'h4b301;
         mem[293] =  20'h45da2;
         mem[294] =  20'h470c3;
         mem[295] =  20'h57a02;
         mem[296] =  20'h624c3;
         mem[297] =  20'h5dcc3;
         mem[298] =  20'h2dca4;
         mem[299] =  20'h2e449;
         mem[300] =  20'h03449;
         mem[301] =  20'h02449;
         mem[302] =  20'h1644f;
         mem[303] =  20'h14c4f;
         mem[304] =  20'h1cd22;
         mem[305] =  20'h40867;
         mem[306] =  20'h790c5;
         mem[307] =  20'h6c0a4;
         mem[308] =  20'h54c68;
         mem[309] =  20'h71241;
         mem[310] =  20'h78261;
         mem[311] =  20'h02c49;
         mem[312] =  20'h1c432;
         mem[313] =  20'h1b832;
         mem[314] =  20'h150c9;
         mem[315] =  20'h0844e;
         mem[316] =  20'h79d23;
         mem[317] =  20'h13148;
         mem[318] =  20'h23066;
         mem[319] =  20'h0cd68;
         mem[320] =  20'h794a5;
         mem[321] =  20'h8a641;
         mem[322] =  20'h5a84a;
         mem[323] =  20'h0e904;
         mem[324] =  20'h2d583;
         mem[325] =  20'h28085;
         mem[326] =  20'h4c5c4;
         mem[327] =  20'h58885;
         mem[328] =  20'h540a7;
         mem[329] =  20'h59468;
         mem[330] =  20'h2e0c8;
         mem[331] =  20'h19a81;
         mem[332] =  20'h58662;
         mem[333] =  20'h28049;
         mem[334] =  20'h2986e;
         mem[335] =  20'h3a84c;
         mem[336] =  20'h2ac69;
         mem[337] =  20'h25869;
         mem[338] =  20'h23cc3;
         mem[339] =  20'h7dde2;
         mem[340] =  20'h23cc3;
         mem[341] =  20'h1f4c3;
         mem[342] =  20'h46241;
         mem[343] =  20'h0e182;
         mem[344] =  20'h03049;
         mem[345] =  20'h02849;
         mem[346] =  20'h5b522;
         mem[347] =  20'h32da2;
         mem[348] =  20'h5b522;
         mem[349] =  20'h2086f;
         mem[350] =  20'h34c66;
         mem[351] =  20'h53467;
         mem[352] =  20'h5b522;
         mem[353] =  20'h4d4a4;
         mem[354] =  20'h09853;
         mem[355] =  20'h08853;
         mem[356] =  20'h4f8c3;
         mem[357] =  20'h89e41;
         mem[358] =  20'h67943;
         mem[359] =  20'h51962;
         mem[360] =  20'h28903;
         mem[361] =  20'h0052b;
         mem[362] =  20'h2f487;
         mem[363] =  20'h1906a;
         mem[364] =  20'h04449;
         mem[365] =  20'h01449;
         mem[366] =  20'h4f866;
         mem[367] =  20'h4bc66;
         mem[368] =  20'h5b522;
         mem[369] =  20'h57922;
         mem[370] =  20'h5ee61;
         mem[371] =  20'h58261;
         mem[372] =  20'h6dd42;
         mem[373] =  20'h018a6;
         mem[374] =  20'h0b466;
         mem[375] =  20'h06866;
         mem[376] =  20'h6e4c3;
         mem[377] =  20'h3a126;
         mem[378] =  20'h2ec86;
         mem[379] =  20'h1a1c4;
         mem[380] =  20'h28849;
         mem[381] =  20'h408c3;
         mem[382] =  20'h6e122;
         mem[383] =  20'h080f7;
         mem[384] =  20'h46622;
         mem[385] =  20'h25d66;
         mem[386] =  20'h6bda2;
         mem[387] =  20'h6a522;
         mem[388] =  20'h2f0a4;
         mem[389] =  20'h600c3;
         mem[390] =  20'h350c3;
         mem[391] =  20'h59904;
         mem[392] =  20'h68066;
         mem[393] =  20'h19301;
         mem[394] =  20'h7a542;
         mem[395] =  20'h530c3;
         mem[396] =  20'h14243;
         mem[397] =  20'h26a03;
         mem[398] =  20'h48c66;
         mem[399] =  20'h2d4c4;
         mem[400] =  20'h28849;
         mem[401] =  20'h34c4a;
         mem[402] =  20'h60849;
         mem[403] =  20'h09535;
         mem[404] =  20'h338c7;
         mem[405] =  20'h21c49;
         mem[406] =  20'h0e904;
         mem[407] =  20'h484a4;
         mem[408] =  20'h460a4;
         mem[409] =  20'h28449;
         mem[410] =  20'h07071;
         mem[411] =  20'h19e63;
         mem[412] =  20'h714c3;
         mem[413] =  20'h1e053;
         mem[414] =  20'h654a7;
         mem[415] =  20'h2f0a6;
         mem[416] =  20'h2d4a6;
         mem[417] =  20'h0f866;
         mem[418] =  20'h7f0e4;
         mem[419] =  20'h59d22;
         mem[420] =  20'h0f066;
         mem[421] =  20'h0344e;
         mem[422] =  20'h0244e;
         mem[423] =  20'h6dd22;
         mem[424] =  20'h340c5;
         mem[425] =  20'h17c4b;
         mem[426] =  20'h4c967;
         mem[427] =  20'h304c3;
         mem[428] =  20'h33d22;
         mem[429] =  20'h304c3;
         mem[430] =  20'h2bcc3;
         mem[431] =  20'h27d22;
         mem[432] =  20'h8fe61;
         mem[433] =  20'h6e8c3;
         mem[434] =  20'h6a8c3;
         mem[435] =  20'h48449;
         mem[436] =  20'h46c49;
         mem[437] =  20'h3a8c7;
         mem[438] =  20'h6c8c5;
         mem[439] =  20'h03849;
         mem[440] =  20'h02049;
         mem[441] =  20'h72241;
         mem[442] =  20'h70e41;
         mem[443] =  20'h4d966;
         mem[444] =  20'h26ce3;
         mem[445] =  20'h26de2;
         mem[446] =  20'h066c1;
         mem[447] =  20'h02118;
         mem[448] =  20'h60524;
         mem[449] =  20'h46583;
         mem[450] =  20'h650e4;
         mem[451] =  20'h0f963;
         mem[452] =  20'h800e3;
         mem[453] =  20'h03188;
         mem[454] =  20'h52122;
         mem[455] =  20'h456c1;
         mem[456] =  20'h2d564;
         mem[457] =  20'h358c3;
         mem[458] =  20'h38702;
         mem[459] =  20'h04ca5;
         mem[460] =  20'h000a5;
         mem[461] =  20'h09582;
         mem[462] =  20'h70a41;
         mem[463] =  20'h61103;
         mem[464] =  20'h5e903;
         mem[465] =  20'h6be41;
         mem[466] =  20'h70aa5;
         mem[467] =  20'h03c58;
         mem[468] =  20'h1b44b;
         mem[469] =  20'h22466;
         mem[470] =  20'h57c4a;
         mem[471] =  20'h03c58;
         mem[472] =  20'h01c58;
         mem[473] =  20'h30867;
         mem[474] =  20'h2d44c;
         mem[475] =  20'h2150e;
         mem[476] =  20'h5f142;
         mem[477] =  20'h03849;
         mem[478] =  20'h2c467;
         mem[479] =  20'h1106f;
         mem[480] =  20'h0d049;
         mem[481] =  20'h10ca7;
         mem[482] =  20'h28832;
         mem[483] =  20'h22ca6;
         mem[484] =  20'h2804a;
         mem[485] =  20'h03849;
         mem[486] =  20'h14467;
         mem[487] =  20'h2d4e3;
         mem[488] =  20'h2e886;
         mem[489] =  20'h544e6;
         mem[490] =  20'h28049;
         mem[491] =  20'h6e4c3;
         mem[492] =  20'h0184d;
         mem[493] =  20'h0ece3;
         mem[494] =  20'h334a4;
         mem[495] =  20'h34885;
         mem[496] =  20'h340a4;
         mem[497] =  20'h14563;
         mem[498] =  20'h28085;
         mem[499] =  20'h02105;
         mem[500] =  20'h4b6e2;
         mem[501] =  20'h858c3;
         mem[502] =  20'h32ea2;
         mem[503] =  20'h1fc4c;
         mem[504] =  20'h2e485;
         mem[505] =  20'h4d105;
         mem[506] =  20'h2e4ac;
         mem[507] =  20'h76d42;
         mem[508] =  20'h80922;
         mem[509] =  20'h59cc8;
         mem[510] =  20'h80922;
         mem[511] =  20'h7d522;
         mem[512] =  20'h48922;
         mem[513] =  20'h44d22;
         mem[514] =  20'h17849;
         mem[515] =  20'h71241;
         mem[516] =  20'h6b2a2;
         mem[517] =  20'h7f4c3;
         mem[518] =  20'h2a0c3;
         mem[519] =  20'h258c3;
         mem[520] =  20'h03105;
         mem[521] =  20'h008a8;
         mem[522] =  20'h038a5;
         mem[523] =  20'h014a5;
         mem[524] =  20'h1746a;
         mem[525] =  20'h460c3;
         mem[526] =  20'h05832;
         mem[527] =  20'h02049;
         mem[528] =  20'h34c67;
         mem[529] =  20'h4cc85;
         mem[530] =  20'h05832;
         mem[531] =  20'h28849;
         mem[532] =  20'h10522;
         mem[533] =  20'h12f01;
         mem[534] =  20'h2f049;
         mem[535] =  20'h27c4a;
         mem[536] =  20'h09c4c;
         mem[537] =  20'h40186;
         mem[538] =  20'h16435;
         mem[539] =  20'h20d84;
         mem[540] =  20'h19e44;
         mem[541] =  20'h07241;
         mem[542] =  20'h54582;
         mem[543] =  20'h22449;
         mem[544] =  20'h09849;
         mem[545] =  20'h0e856;
         mem[546] =  20'h43887;
         mem[547] =  20'h39205;
         mem[548] =  20'h43887;
         mem[549] =  20'h3e887;
         mem[550] =  20'h6cd63;
         mem[551] =  20'h2dd09;
         mem[552] =  20'h09850;
         mem[553] =  20'h08850;
         mem[554] =  20'h22904;
         mem[555] =  20'h4b0c3;
         mem[556] =  20'h6be41;
         mem[557] =  20'h5e8c3;
         mem[558] =  20'h66122;
         mem[559] =  20'h51c85;
         mem[560] =  20'h48866;
         mem[561] =  20'h26641;
         mem[562] =  20'h2404b;
         mem[563] =  20'h2004b;
         mem[564] =  20'h0b049;
         mem[565] =  20'h07049;
         mem[566] =  20'h5ed29;
         mem[567] =  20'h46582;
         mem[568] =  20'h1cd22;
         mem[569] =  20'h19122;
         mem[570] =  20'h04451;
         mem[571] =  20'h01451;
         mem[572] =  20'h78d22;
         mem[573] =  20'h46466;
         mem[574] =  20'h335c6;
         mem[575] =  20'h34866;
         mem[576] =  20'h4d9c5;
         mem[577] =  20'h4b1c5;
         mem[578] =  20'h10522;
         mem[579] =  20'h0c922;
         mem[580] =  20'h2904e;
         mem[581] =  20'h2e849;
         mem[582] =  20'h2904f;
         mem[583] =  20'h2784f;
         mem[584] =  20'h16889;
         mem[585] =  20'h00c75;
         mem[586] =  20'h54104;
         mem[587] =  20'h2d4a6;
         mem[588] =  20'h28849;
         mem[589] =  20'h12cc3;
         mem[590] =  20'h5ea41;
         mem[591] =  20'h58485;
         mem[592] =  20'h4e182;
         mem[593] =  20'h0cc34;
         mem[594] =  20'h684a4;
         mem[595] =  20'h648a4;
         mem[596] =  20'h14943;
         mem[597] =  20'h02103;
         mem[598] =  20'h3f5e2;
         mem[599] =  20'h21c86;
         mem[600] =  20'h655c3;
         mem[601] =  20'h79885;
         mem[602] =  20'h26467;
         mem[603] =  20'h04866;
         mem[604] =  20'h0d641;
         mem[605] =  20'h4d5c6;
         mem[606] =  20'h00c66;
         mem[607] =  20'h48066;
         mem[608] =  20'h7f103;
         mem[609] =  20'h48067;
         mem[610] =  20'h58942;
         mem[611] =  20'h48066;
         mem[612] =  20'h46c67;
         mem[613] =  20'h33d64;
         mem[614] =  20'h6bd42;
         mem[615] =  20'h04049;
         mem[616] =  20'h01849;
         mem[617] =  20'h2e885;
         mem[618] =  20'h06681;
         mem[619] =  20'h80542;
         mem[620] =  20'h2d06b;
         mem[621] =  20'h6cd43;
         mem[622] =  20'h0f049;
         mem[623] =  20'h164a4;
         mem[624] =  20'h270c3;
         mem[625] =  20'h35085;
         mem[626] =  20'h4cc88;
         mem[627] =  20'h40922;
         mem[628] =  20'h209c3;
         mem[629] =  20'h7de64;
         mem[630] =  20'h014a8;
         mem[631] =  20'h0dd12;
         mem[632] =  20'h46d0b;
         mem[633] =  20'h13925;
         mem[634] =  20'h6aa41;
         mem[635] =  20'h71e41;
         mem[636] =  20'h5e122;
         mem[637] =  20'h57ee5;
         mem[638] =  20'h32e41;
         mem[639] =  20'h338c3;
         mem[640] =  20'h0e436;
         mem[641] =  20'h7a542;
         mem[642] =  20'h7d542;
         mem[643] =  20'h1604c;
         mem[644] =  20'h28849;
         mem[645] =  20'h03449;
         mem[646] =  20'h02449;
         mem[647] =  20'h42466;
         mem[648] =  20'h46069;
         mem[649] =  20'h23033;
         mem[650] =  20'h33922;
         mem[651] =  20'h23033;
         mem[652] =  20'h258c3;
         mem[653] =  20'h8ae41;
         mem[654] =  20'h404c4;
         mem[655] =  20'h1d485;
         mem[656] =  20'h34866;
         mem[657] =  20'h3c068;
         mem[658] =  20'h3e8a4;
         mem[659] =  20'h290e3;
         mem[660] =  20'h21433;
         mem[661] =  20'h1c4b4;
         mem[662] =  20'h1a8b4;
         mem[663] =  20'h41c66;
         mem[664] =  20'h40866;
         mem[665] =  20'h10c67;
         mem[666] =  20'h0d867;
         mem[667] =  20'h1c067;
         mem[668] =  20'h1bc49;
         mem[669] =  20'h1bc8a;
         mem[670] =  20'h1b48a;
         mem[671] =  20'h7f142;
         mem[672] =  20'h7d6a2;
         mem[673] =  20'h0ecc6;
         mem[674] =  20'h0ecc6;
         mem[675] =  20'h23cc3;
         mem[676] =  20'h46cc3;
         mem[677] =  20'h38e82;
         mem[678] =  20'h1f4c3;
         mem[679] =  20'h5c085;
         mem[680] =  20'h58085;
         mem[681] =  20'h4554d;
         mem[682] =  20'h3b4c5;
         mem[683] =  20'h28d03;
         mem[684] =  20'h83922;
         mem[685] =  20'h22085;
         mem[686] =  20'h200e6;
         mem[687] =  20'h1c066;
         mem[688] =  20'h2c661;
         mem[689] =  20'h55cc3;
         mem[690] =  20'h32e41;
         mem[691] =  20'h12049;
         mem[692] =  20'h77681;
         mem[693] =  20'h3eec1;
         mem[694] =  20'h0c849;
         mem[695] =  20'h04c57;
         mem[696] =  20'h13873;
         mem[697] =  20'h11849;
         mem[698] =  20'h2bd42;
         mem[699] =  20'h034c6;
         mem[700] =  20'h12d83;
         mem[701] =  20'h79485;
         mem[702] =  20'h59885;
         mem[703] =  20'h58a23;
         mem[704] =  20'h1fd24;
         mem[705] =  20'h290e3;
         mem[706] =  20'h264e3;
         mem[707] =  20'h23832;
         mem[708] =  20'h20c32;
         mem[709] =  20'h4d9c2;
         mem[710] =  20'h4c122;
         mem[711] =  20'h13643;
         mem[712] =  20'h15488;
         mem[713] =  20'h07885;
         mem[714] =  20'h47ce4;
         mem[715] =  20'h57ac2;
         mem[716] =  20'h48885;
         mem[717] =  20'h460e4;
         mem[718] =  20'h7f122;
         mem[719] =  20'h196c2;
         mem[720] =  20'h17851;
         mem[721] =  20'h46d09;
         mem[722] =  20'h05066;
         mem[723] =  20'h02449;
         mem[724] =  20'h48926;
         mem[725] =  20'h90641;
         mem[726] =  20'h428c3;
         mem[727] =  20'h06c4b;
         mem[728] =  20'h0504a;
         mem[729] =  20'h13851;
         mem[730] =  20'h6e122;
         mem[731] =  20'h64103;
         mem[732] =  20'h4f0c4;
         mem[733] =  20'h4b8c4;
         mem[734] =  20'h2e485;
         mem[735] =  20'h25e61;
         mem[736] =  20'h35867;
         mem[737] =  20'h45983;
         mem[738] =  20'h2ca41;
         mem[739] =  20'h28086;
         mem[740] =  20'h3912e;
         mem[741] =  20'h00849;
         mem[742] =  20'h22452;
         mem[743] =  20'h21c52;
         mem[744] =  20'h2244a;
         mem[745] =  20'h1bc4b;
         mem[746] =  20'h6b641;
         mem[747] =  20'h6a681;
         mem[748] =  20'h538c4;
         mem[749] =  20'h6c504;
         mem[750] =  20'h67466;
         mem[751] =  20'h398e7;
         mem[752] =  20'h03185;
         mem[753] =  20'h4b641;
         mem[754] =  20'h3d0a4;
         mem[755] =  20'h384a4;
         mem[756] =  20'h2a889;
         mem[757] =  20'h25889;
         mem[758] =  20'h23cc6;
         mem[759] =  20'h27c49;
         mem[760] =  20'h5404b;
         mem[761] =  20'h1f4c6;
         mem[762] =  20'h132e1;
         mem[763] =  20'h64661;
         mem[764] =  20'h7a162;
         mem[765] =  20'h52485;
         mem[766] =  20'h418a4;
         mem[767] =  20'h39523;
         mem[768] =  20'h67d22;
         mem[769] =  20'h57d22;
         mem[770] =  20'h41d44;
         mem[771] =  20'h01472;
         mem[772] =  20'h48c6a;
         mem[773] =  20'h0dc85;
         mem[774] =  20'h1b8e6;
         mem[775] =  20'h01ca7;
         mem[776] =  20'h79d82;
         mem[777] =  20'h322e2;
         mem[778] =  20'h42c85;
         mem[779] =  20'h6a641;
         mem[780] =  20'h74522;
         mem[781] =  20'h70922;
         mem[782] =  20'h48066;
         mem[783] =  20'h46c66;
         mem[784] =  20'h15d83;
         mem[785] =  20'h1fe41;
         mem[786] =  20'h03182;
         mem[787] =  20'h6aa41;
         mem[788] =  20'h6e122;
         mem[789] =  20'h6a522;
         mem[790] =  20'h72241;
         mem[791] =  20'h3484a;
         mem[792] =  20'h28849;
         mem[793] =  20'h4d0a4;
         mem[794] =  20'h4e0c4;
         mem[795] =  20'h2144b;
         mem[796] =  20'h3b903;
         mem[797] =  20'h38aa2;
         mem[798] =  20'h48866;
         mem[799] =  20'h52d64;
         mem[800] =  20'h368a4;
         mem[801] =  20'h34cc3;
         mem[802] =  20'h47cc4;
         mem[803] =  20'h44ecb;
         mem[804] =  20'h284c4;
         mem[805] =  20'h02c49;
         mem[806] =  20'h03049;
         mem[807] =  20'h14c67;
         mem[808] =  20'h40cc8;
         mem[809] =  20'h2e467;
         mem[810] =  20'h5260a;
         mem[811] =  20'h1bc4a;
         mem[812] =  20'h0de02;
         mem[813] =  20'h214c4;
         mem[814] =  20'h03c49;
         mem[815] =  20'h1c085;
         mem[816] =  20'h418a4;
         mem[817] =  20'h404a4;
         mem[818] =  20'h47885;
         mem[819] =  20'h3f485;
         mem[820] =  20'h4e868;
         mem[821] =  20'h85503;
         mem[822] =  20'h7f4c4;
         mem[823] =  20'h6a922;
         mem[824] =  20'h79942;
         mem[825] =  20'h72c86;
         mem[826] =  20'h28866;
         mem[827] =  20'h644c3;
         mem[828] =  20'h72182;
         mem[829] =  20'h25e81;
         mem[830] =  20'h1b123;
         mem[831] =  20'h83d22;
         mem[832] =  20'h2e886;
         mem[833] =  20'h0e486;
         mem[834] =  20'h42068;
         mem[835] =  20'h47085;
         mem[836] =  20'h3bc66;
         mem[837] =  20'h40449;
         mem[838] =  20'h45ca4;
         mem[839] =  20'h024e6;
         mem[840] =  20'h33d42;
         mem[841] =  20'h02c4f;
         mem[842] =  20'h13641;
         mem[843] =  20'h7f103;
         mem[844] =  20'h07241;
         mem[845] =  20'h02c66;
         mem[846] =  20'h70a41;
         mem[847] =  20'h2e485;
         mem[848] =  20'h13449;
         mem[849] =  20'h11849;
         mem[850] =  20'h0d049;
         mem[851] =  20'h09582;
         mem[852] =  20'h70922;
         mem[853] =  20'h61522;
         mem[854] =  20'h64261;
         mem[855] =  20'h22566;
         mem[856] =  20'h53466;
         mem[857] =  20'h13e81;
         mem[858] =  20'h5a04a;
         mem[859] =  20'h4e903;
         mem[860] =  20'h64903;
         mem[861] =  20'h35867;
         mem[862] =  20'h4b903;
         mem[863] =  20'h7e604;
         mem[864] =  20'h2e086;
         mem[865] =  20'h0f885;
         mem[866] =  20'h270c3;
         mem[867] =  20'h2ec49;
         mem[868] =  20'h00086;
         mem[869] =  20'h494c3;
         mem[870] =  20'h4c466;
         mem[871] =  20'h85ce3;
         mem[872] =  20'h13603;
         mem[873] =  20'h3b8e3;
         mem[874] =  20'h46487;
         mem[875] =  20'h2e849;
         mem[876] =  20'h33c67;
         mem[877] =  20'h68888;
         mem[878] =  20'h5a44a;
         mem[879] =  20'h47485;
         mem[880] =  20'h516e1;
         mem[881] =  20'h03c4c;
         mem[882] =  20'h3f885;
         mem[883] =  20'h1c542;
         mem[884] =  20'h01c4c;
         mem[885] =  20'h29066;
         mem[886] =  20'h27466;
         mem[887] =  20'h47ccd;
         mem[888] =  20'h464cd;
         mem[889] =  20'h68086;
         mem[890] =  20'h2bea1;
         mem[891] =  20'h68086;
         mem[892] =  20'h58cc7;
         mem[893] =  20'h46261;
         mem[894] =  20'h26dc2;
         mem[895] =  20'h72cc4;
         mem[896] =  20'h02449;
         mem[897] =  20'h22962;
         mem[898] =  20'h01466;
         mem[899] =  20'h0b057;
         mem[900] =  20'h07057;
         mem[901] =  20'h6ba41;
         mem[902] =  20'h1f562;
         mem[903] =  20'h6ae81;
         mem[904] =  20'h209a2;
         mem[905] =  20'h3896f;
         mem[906] =  20'h1b8e3;
         mem[907] =  20'h2dca4;
         mem[908] =  20'h2e8a4;
         mem[909] =  20'h1c049;
         mem[910] =  20'h4c066;
         mem[911] =  20'h15c85;
         mem[912] =  20'h26503;
         mem[913] =  20'h399c3;
         mem[914] =  20'h20522;
         mem[915] =  20'h1aa41;
         mem[916] =  20'h28066;
         mem[917] =  20'h0cb01;
         mem[918] =  20'h76d42;
         mem[919] =  20'h77a41;
         mem[920] =  20'h1fc68;
         mem[921] =  20'h33d62;
         mem[922] =  20'h5298b;
         mem[923] =  20'h4d885;
         mem[924] =  20'h27c86;
         mem[925] =  20'h494c3;
         mem[926] =  20'h2e0aa;
         mem[927] =  20'h22449;
         mem[928] =  20'h3b04a;
         mem[929] =  20'h5ac4a;
         mem[930] =  20'h59c4a;
         mem[931] =  20'h45e03;
         mem[932] =  20'h4ba81;
         mem[933] =  20'h0344d;
         mem[934] =  20'h0244d;
         mem[935] =  20'h088c7;
         mem[936] =  20'h57cc3;
         mem[937] =  20'h7f122;
         mem[938] =  20'h459e2;
         mem[939] =  20'h46261;
         mem[940] =  20'h598e8;
         mem[941] =  20'h66522;
         mem[942] =  20'h44d04;
         mem[943] =  20'h20e41;
         mem[944] =  20'h65086;
         mem[945] =  20'h61122;
         mem[946] =  20'h334e7;
         mem[947] =  20'h67163;
         mem[948] =  20'h02c49;
         mem[949] =  20'h22ca5;
         mem[950] =  20'h208a5;
         mem[951] =  20'h28903;
         mem[952] =  20'h3e8c3;
         mem[953] =  20'h43887;
         mem[954] =  20'h72cc6;
         mem[955] =  20'h41886;
         mem[956] =  20'h02849;
         mem[957] =  20'h1c888;
         mem[958] =  20'h4cd42;
         mem[959] =  20'h288e7;
         mem[960] =  20'h4ba81;
         mem[961] =  20'h68888;
         mem[962] =  20'h450c5;
         mem[963] =  20'h46582;
         mem[964] =  20'h4e067;
         mem[965] =  20'h1c888;
         mem[966] =  20'h1a888;
         mem[967] =  20'h3b066;
         mem[968] =  20'h1f906;
         mem[969] =  20'h3a868;
         mem[970] =  20'h01c32;
         mem[971] =  20'h684a7;
         mem[972] =  20'h648a7;
         mem[973] =  20'h2d943;
         mem[974] =  20'h38ae6;
         mem[975] =  20'h084e3;
         mem[976] =  20'h28449;
         mem[977] =  20'h714c3;
         mem[978] =  20'h37088;
         mem[979] =  20'h78d04;
         mem[980] =  20'h37088;
         mem[981] =  20'h32088;
         mem[982] =  20'h6c505;
         mem[983] =  20'h460a4;
         mem[984] =  20'h0da61;
         mem[985] =  20'h4d109;
         mem[986] =  20'h1a9a4;
         mem[987] =  20'h06701;
         mem[988] =  20'h17c4b;
         mem[989] =  20'h28049;
         mem[990] =  20'h47cc4;
         mem[991] =  20'h320c3;
         mem[992] =  20'h72241;
         mem[993] =  20'h64122;
         mem[994] =  20'h17c49;
         mem[995] =  20'h13449;
         mem[996] =  20'h04873;
         mem[997] =  20'h00c73;
         mem[998] =  20'h48068;
         mem[999] =  20'h46c68;
         mem[1000] =  20'h4c661;
         mem[1001] =  20'h7f4c4;
         mem[1002] =  20'h33a02;
         mem[1003] =  20'h02466;
         mem[1004] =  20'h41087;
         mem[1005] =  20'h451e6;
         mem[1006] =  20'h4dc85;
         mem[1007] =  20'h01c49;
         mem[1008] =  20'h03849;
         mem[1009] =  20'h208c4;
         mem[1010] =  20'h5ad62;
         mem[1011] =  20'h57aa1;
         mem[1012] =  20'h09486;
         mem[1013] =  20'h00466;
         mem[1014] =  20'h136a1;
         mem[1015] =  20'h13661;
         mem[1016] =  20'h43867;
         mem[1017] =  20'h3ec67;
         mem[1018] =  20'h290e7;
         mem[1019] =  20'h57922;
         mem[1020] =  20'h6e103;
         mem[1021] =  20'h06962;
         mem[1022] =  20'h53922;
         mem[1023] =  20'h64241;
         mem[1024] =  20'h6e4e3;
         mem[1025] =  20'h15d04;
         mem[1026] =  20'h274c5;
         mem[1027] =  20'h28449;
         mem[1028] =  20'h0944a;
         mem[1029] =  20'h08c4a;
         mem[1030] =  20'h744c3;
         mem[1031] =  20'h714c3;
         mem[1032] =  20'h0a433;
         mem[1033] =  20'h13849;
         mem[1034] =  20'h04033;
         mem[1035] =  20'h15cc4;
         mem[1036] =  20'h21c49;
         mem[1037] =  20'h01c33;
         mem[1038] =  20'h2e866;
         mem[1039] =  20'h2e8a5;
         mem[1040] =  20'h15c32;
         mem[1041] =  20'h1584c;
         mem[1042] =  20'h32e61;
         mem[1043] =  20'h32a41;
         mem[1044] =  20'h54522;
         mem[1045] =  20'h20849;
         mem[1046] =  20'h09d42;
         mem[1047] =  20'h06542;
         mem[1048] =  20'h60466;
         mem[1049] =  20'h0e908;
         mem[1050] =  20'h26e41;
         mem[1051] =  20'h60866;
         mem[1052] =  20'h4dc85;
         mem[1053] =  20'h4d485;
         mem[1054] =  20'h0ddc2;
         mem[1055] =  20'h2e485;
         mem[1056] =  20'h474a4;
         mem[1057] =  20'h3a087;
         mem[1058] =  20'h22563;
         mem[1059] =  20'h320c3;
         mem[1060] =  20'h79d22;
         mem[1061] =  20'h77661;
         mem[1062] =  20'h79d22;
         mem[1063] =  20'h70e41;
         mem[1064] =  20'h79d22;
         mem[1065] =  20'h06701;
         mem[1066] =  20'h0ddc2;
         mem[1067] =  20'h65922;
         mem[1068] =  20'h678c3;
         mem[1069] =  20'h8ada2;
         mem[1070] =  20'h538c4;
         mem[1071] =  20'h408e3;
         mem[1072] =  20'h34c66;
         mem[1073] =  20'h40067;
         mem[1074] =  20'h42ca4;
         mem[1075] =  20'h5fd03;
         mem[1076] =  20'h2dd22;
         mem[1077] =  20'h650c3;
         mem[1078] =  20'h79d22;
         mem[1079] =  20'h600c3;
         mem[1080] =  20'h3c4e5;
         mem[1081] =  20'h388e5;
         mem[1082] =  20'h2e871;
         mem[1083] =  20'h19c6a;
         mem[1084] =  20'h33ca4;
         mem[1085] =  20'h2ec49;
         mem[1086] =  20'h60c49;
         mem[1087] =  20'h32c68;
         mem[1088] =  20'h79d22;
         mem[1089] =  20'h77922;
         mem[1090] =  20'h09866;
         mem[1091] =  20'h4c485;
         mem[1092] =  20'h22086;
         mem[1093] =  20'h1b468;
         mem[1094] =  20'h684a4;
         mem[1095] =  20'h648a4;
         mem[1096] =  20'h03182;
         mem[1097] =  20'h32122;
         mem[1098] =  20'h1c183;
         mem[1099] =  20'h0dd62;
         mem[1100] =  20'h09562;
         mem[1101] =  20'h600c9;
         mem[1102] =  20'h45682;
         mem[1103] =  20'h399c7;
         mem[1104] =  20'h20603;
         mem[1105] =  20'h19a61;
         mem[1106] =  20'h14942;
         mem[1107] =  20'h57885;
         mem[1108] =  20'h456a1;
         mem[1109] =  20'h01866;
         mem[1110] =  20'h2d5c3;
         mem[1111] =  20'h09049;
         mem[1112] =  20'h48923;
         mem[1113] =  20'h2dc87;
         mem[1114] =  20'h90a61;
         mem[1115] =  20'h64a81;
         mem[1116] =  20'h04c4d;
         mem[1117] =  20'h45104;
         mem[1118] =  20'h6dcc3;
         mem[1119] =  20'h6b4c3;
         mem[1120] =  20'h22c4a;
         mem[1121] =  20'h2144a;
         mem[1122] =  20'h358c3;
         mem[1123] =  20'h330c3;
         mem[1124] =  20'h0e915;
         mem[1125] =  20'h0d44d;
         mem[1126] =  20'h05055;
         mem[1127] =  20'h19854;
         mem[1128] =  20'h72922;
         mem[1129] =  20'h02449;
         mem[1130] =  20'h61ce3;
         mem[1131] =  20'h864e3;
         mem[1132] =  20'h22069;
         mem[1133] =  20'h2244a;
         mem[1134] =  20'h28849;
         mem[1135] =  20'h21c69;
         mem[1136] =  20'h67942;
         mem[1137] =  20'h208e7;
         mem[1138] =  20'h368c3;
         mem[1139] =  20'h270c6;
         mem[1140] =  20'h5484a;
         mem[1141] =  20'h3ed44;
         mem[1142] =  20'h61922;
         mem[1143] =  20'h150c3;
         mem[1144] =  20'h348a7;
         mem[1145] =  20'h26602;
         mem[1146] =  20'h29903;
         mem[1147] =  20'h5384a;
         mem[1148] =  20'h61922;
         mem[1149] =  20'h5dd22;
         mem[1150] =  20'h73d22;
         mem[1151] =  20'h71122;
         mem[1152] =  20'h6ba41;
         mem[1153] =  20'h6aa41;
         mem[1154] =  20'h07a41;
         mem[1155] =  20'h0ce61;
         mem[1156] =  20'h1084b;
         mem[1157] =  20'h600a6;
         mem[1158] =  20'h1084b;
         mem[1159] =  20'h0e04b;
         mem[1160] =  20'h23cc3;
         mem[1161] =  20'h0cd62;
         mem[1162] =  20'h024ec;
         mem[1163] =  20'h51641;
         mem[1164] =  20'h10049;
         mem[1165] =  20'h45a41;
         mem[1166] =  20'h29903;
         mem[1167] =  20'h32e41;
         mem[1168] =  20'h47849;
         mem[1169] =  20'h34c49;
         mem[1170] =  20'h03c32;
         mem[1171] =  20'h02032;
         mem[1172] =  20'h29ce3;
         mem[1173] =  20'h7dd22;
         mem[1174] =  20'h77aa1;
         mem[1175] =  20'h258e3;
         mem[1176] =  20'h32ac1;
         mem[1177] =  20'h12d88;
         mem[1178] =  20'h7a122;
         mem[1179] =  20'h208c4;
         mem[1180] =  20'h288e3;
         mem[1181] =  20'h654e3;
         mem[1182] =  20'h23cc3;
         mem[1183] =  20'h1f4c3;
         mem[1184] =  20'h1c545;
         mem[1185] =  20'h52868;
         mem[1186] =  20'h088ef;
         mem[1187] =  20'h4e0e8;
         mem[1188] =  20'h2d4c4;
         mem[1189] =  20'h21866;
         mem[1190] =  20'h48066;
         mem[1191] =  20'h46c66;
         mem[1192] =  20'h20e41;
         mem[1193] =  20'h0d04b;
         mem[1194] =  20'h0504f;
         mem[1195] =  20'h0084d;
         mem[1196] =  20'h03849;
         mem[1197] =  20'h02049;
         mem[1198] =  20'h0e904;
         mem[1199] =  20'h54524;
         mem[1200] =  20'h2e0a4;
         mem[1201] =  20'h34cc3;
         mem[1202] =  20'h5ee61;
         mem[1203] =  20'h4108a;
         mem[1204] =  20'h6c522;
         mem[1205] =  20'h3a0a4;
         mem[1206] =  20'h1c087;
         mem[1207] =  20'h514c3;
         mem[1208] =  20'h368c3;
         mem[1209] =  20'h70903;
         mem[1210] =  20'h748e3;
         mem[1211] =  20'h7d542;
         mem[1212] =  20'h35143;
         mem[1213] =  20'h34449;
         mem[1214] =  20'h22488;
         mem[1215] =  20'h21488;
         mem[1216] =  20'h28849;
         mem[1217] =  20'h01050;
         mem[1218] =  20'h35cc4;
         mem[1219] =  20'h32cc4;
         mem[1220] =  20'h5b522;
         mem[1221] =  20'h45deb;
         mem[1222] =  20'h5b522;
         mem[1223] =  20'h57922;
         mem[1224] =  20'h6e122;
         mem[1225] =  20'h6a522;
         mem[1226] =  20'h03885;
         mem[1227] =  20'h00c50;
         mem[1228] =  20'h33d42;
         mem[1229] =  20'h6cc85;
         mem[1230] =  20'h27942;
         mem[1231] =  20'h8c922;
         mem[1232] =  20'h3a162;
         mem[1233] =  20'h000c5;
         mem[1234] =  20'h0a4c3;
         mem[1235] =  20'h72522;
         mem[1236] =  20'h2e4b0;
         mem[1237] =  20'h414cd;
         mem[1238] =  20'h0f8c3;
         mem[1239] =  20'h4bd83;
         mem[1240] =  20'h23503;
         mem[1241] =  20'h1f503;
         mem[1242] =  20'h12d8b;
         mem[1243] =  20'h51485;
         mem[1244] =  20'h79485;
         mem[1245] =  20'h3ac87;
         mem[1246] =  20'h2cde3;
         mem[1247] =  20'h08506;
         mem[1248] =  20'h59ca8;
         mem[1249] =  20'h858c3;
         mem[1250] =  20'h46466;
         mem[1251] =  20'h28449;
         mem[1252] =  20'h27868;
         mem[1253] =  20'h1a281;
         mem[1254] =  20'h408c3;
         mem[1255] =  20'h6c142;
         mem[1256] =  20'h19449;
         mem[1257] =  20'h03c49;
         mem[1258] =  20'h01c49;
         mem[1259] =  20'h03449;
         mem[1260] =  20'h2e066;
         mem[1261] =  20'h07241;
         mem[1262] =  20'h3e942;
         mem[1263] =  20'h34886;
         mem[1264] =  20'h20c66;
         mem[1265] =  20'h03d2b;
         mem[1266] =  20'h0012b;
         mem[1267] =  20'h1184b;
         mem[1268] =  20'h0d04b;
         mem[1269] =  20'h03449;
         mem[1270] =  20'h06681;
         mem[1271] =  20'h13681;
         mem[1272] =  20'h45241;
         mem[1273] =  20'h430c3;
         mem[1274] =  20'h12ec3;
         mem[1275] =  20'h29cc3;
         mem[1276] =  20'h3e8c3;
         mem[1277] =  20'h32302;
         mem[1278] =  20'h0d04a;
         mem[1279] =  20'h28849;
         mem[1280] =  20'h02449;
         mem[1281] =  20'h04449;
         mem[1282] =  20'h01449;
         mem[1283] =  20'h7a922;
         mem[1284] =  20'h70a41;
         mem[1285] =  20'h67d22;
         mem[1286] =  20'h6a6e2;
         mem[1287] =  20'h65641;
         mem[1288] =  20'h64122;
         mem[1289] =  20'h35485;
         mem[1290] =  20'h2dca6;
         mem[1291] =  20'h35485;
         mem[1292] =  20'h0206c;
         mem[1293] =  20'h35485;
         mem[1294] =  20'h21c49;
         mem[1295] =  20'h28849;
         mem[1296] =  20'h2e8c4;
         mem[1297] =  20'h35485;
         mem[1298] =  20'h33c85;
         mem[1299] =  20'h42067;
         mem[1300] =  20'h22473;
         mem[1301] =  20'h4e0c3;
         mem[1302] =  20'h38923;
         mem[1303] =  20'h5c885;
         mem[1304] =  20'h38564;
         mem[1305] =  20'h740c3;
         mem[1306] =  20'h25949;
         mem[1307] =  20'h28d46;
         mem[1308] =  20'h640a4;
         mem[1309] =  20'h6be41;
         mem[1310] =  20'h4b261;
         mem[1311] =  20'h3bcc3;
         mem[1312] =  20'h2c162;
         mem[1313] =  20'h41ce4;
         mem[1314] =  20'h3f963;
         mem[1315] =  20'h42ca4;
         mem[1316] =  20'h4c467;
         mem[1317] =  20'h6e4c3;
         mem[1318] =  20'h64cc4;
         mem[1319] =  20'h678c3;
         mem[1320] =  20'h02849;
         mem[1321] =  20'h09057;
         mem[1322] =  20'h70922;
         mem[1323] =  20'h71a41;
         mem[1324] =  20'h399a7;
         mem[1325] =  20'h04c86;
         mem[1326] =  20'h00086;
         mem[1327] =  20'h0e887;
         mem[1328] =  20'h07049;
         mem[1329] =  20'h36466;
         mem[1330] =  20'h33066;
         mem[1331] =  20'h428a5;
         mem[1332] =  20'h3f4a5;
         mem[1333] =  20'h304c3;
         mem[1334] =  20'h4b4c5;
         mem[1335] =  20'h620c4;
         mem[1336] =  20'h0c982;
         mem[1337] =  20'h0a033;
         mem[1338] =  20'h08433;
         mem[1339] =  20'h0bc34;
         mem[1340] =  20'h06834;
         mem[1341] =  20'h49c4c;
         mem[1342] =  20'h4544c;
         mem[1343] =  20'h52247;
         mem[1344] =  20'h590e4;
         mem[1345] =  20'h53184;
         mem[1346] =  20'h73525;
         mem[1347] =  20'h8aa81;
         mem[1348] =  20'h4d466;
         mem[1349] =  20'h2ce41;
         mem[1350] =  20'h2ca41;
         mem[1351] =  20'h304c3;
         mem[1352] =  20'h58122;
         mem[1353] =  20'h5ad22;
         mem[1354] =  20'h2d867;
         mem[1355] =  20'h548c3;
         mem[1356] =  20'h2e489;
         mem[1357] =  20'h4e066;
         mem[1358] =  20'h2bc85;
         mem[1359] =  20'h02c66;
         mem[1360] =  20'h4b983;
         mem[1361] =  20'h548c3;
         mem[1362] =  20'h528c3;
         mem[1363] =  20'h6c922;
         mem[1364] =  20'h78183;
         mem[1365] =  20'h13a81;
         mem[1366] =  20'h20c86;
         mem[1367] =  20'h03038;
         mem[1368] =  20'h660a4;
         mem[1369] =  20'h72cc6;
         mem[1370] =  20'h5e0c4;
         mem[1371] =  20'h43487;
         mem[1372] =  20'h38887;
         mem[1373] =  20'h66525;
         mem[1374] =  20'h39d82;
         mem[1375] =  20'h60c49;
         mem[1376] =  20'h34867;
         mem[1377] =  20'h1c885;
         mem[1378] =  20'h394c3;
         mem[1379] =  20'h2790c;
         mem[1380] =  20'h2d46e;
         mem[1381] =  20'h4fca4;
         mem[1382] =  20'h4b0a4;
         mem[1383] =  20'h29cc3;
         mem[1384] =  20'h25cc3;
         mem[1385] =  20'h23cc3;
         mem[1386] =  20'h1f4c3;
         mem[1387] =  20'h20242;
         mem[1388] =  20'h1fd22;
         mem[1389] =  20'h164a4;
         mem[1390] =  20'h140a4;
         mem[1391] =  20'h4746c;
         mem[1392] =  20'h4786b;
         mem[1393] =  20'h33ca4;
         mem[1394] =  20'h28867;
         mem[1395] =  20'h78241;
         mem[1396] =  20'h1b849;
         mem[1397] =  20'h09067;
         mem[1398] =  20'h47066;
         mem[1399] =  20'h4e84b;
         mem[1400] =  20'h4d04b;
         mem[1401] =  20'h03092;
         mem[1402] =  20'h4cca5;
         mem[1403] =  20'h83ec1;
         mem[1404] =  20'h19434;
         mem[1405] =  20'h0e904;
         mem[1406] =  20'h40542;
         mem[1407] =  20'h2d485;
         mem[1408] =  20'h04467;
         mem[1409] =  20'h5eca4;
         mem[1410] =  20'h13683;
         mem[1411] =  20'h2d4c4;
         mem[1412] =  20'h7f4c3;
         mem[1413] =  20'h4cd42;
         mem[1414] =  20'h21c89;
         mem[1415] =  20'h46c68;
         mem[1416] =  20'h1d851;
         mem[1417] =  20'h00c66;
         mem[1418] =  20'h1d851;
         mem[1419] =  20'h1a051;
         mem[1420] =  20'h78261;
         mem[1421] =  20'h3b049;
         mem[1422] =  20'h55049;
         mem[1423] =  20'h53049;
         mem[1424] =  20'h47ca4;
         mem[1425] =  20'h28849;
         mem[1426] =  20'h03049;
         mem[1427] =  20'h38d04;
         mem[1428] =  20'h740c3;
         mem[1429] =  20'h2e449;
         mem[1430] =  20'h740c3;
         mem[1431] =  20'h58582;
         mem[1432] =  20'h5b122;
         mem[1433] =  20'h57d22;
         mem[1434] =  20'h32e41;
         mem[1435] =  20'h38ac2;
         mem[1436] =  20'h304c3;
         mem[1437] =  20'h2bcc3;
         mem[1438] =  20'h58e03;
         mem[1439] =  20'h72122;
         mem[1440] =  20'h740c3;
         mem[1441] =  20'h718c3;
         mem[1442] =  20'h0a857;
         mem[1443] =  20'h85503;
         mem[1444] =  20'h7f104;
         mem[1445] =  20'h07857;
         mem[1446] =  20'h71641;
         mem[1447] =  20'h6a641;
         mem[1448] =  20'h67162;
         mem[1449] =  20'h70922;
         mem[1450] =  20'h40ce3;
         mem[1451] =  20'h710c3;
         mem[1452] =  20'h2bf02;
         mem[1453] =  20'h2e485;
         mem[1454] =  20'h53cc6;
         mem[1455] =  20'h27849;
         mem[1456] =  20'h03449;
         mem[1457] =  20'h2e849;
         mem[1458] =  20'h0d281;
         mem[1459] =  20'h70cc3;
         mem[1460] =  20'h0fc4d;
         mem[1461] =  20'h2ecc4;
         mem[1462] =  20'h08c4d;
         mem[1463] =  20'h01c32;
         mem[1464] =  20'h164a5;
         mem[1465] =  20'h60488;
         mem[1466] =  20'h41449;
         mem[1467] =  20'h15449;
         mem[1468] =  20'h05067;
         mem[1469] =  20'h00467;
         mem[1470] =  20'h04468;
         mem[1471] =  20'h1b44a;
         mem[1472] =  20'h6d523;
         mem[1473] =  20'h80164;
         mem[1474] =  20'h164a5;
         mem[1475] =  20'h140a5;
         mem[1476] =  20'h29890;
         mem[1477] =  20'h26890;
         mem[1478] =  20'h5a0a5;
         mem[1479] =  20'h772a1;
         mem[1480] =  20'h10522;
         mem[1481] =  20'h094c4;
         mem[1482] =  20'h030c6;
         mem[1483] =  20'h40886;
         mem[1484] =  20'h68ca4;
         mem[1485] =  20'h640a4;
         mem[1486] =  20'h4e885;
         mem[1487] =  20'h658a4;
         mem[1488] =  20'h28cc3;
         mem[1489] =  20'h27c49;
         mem[1490] =  20'h3b867;
         mem[1491] =  20'h3a467;
         mem[1492] =  20'h40566;
         mem[1493] =  20'h33068;
         mem[1494] =  20'h42c87;
         mem[1495] =  20'h3f487;
         mem[1496] =  20'h09c89;
         mem[1497] =  20'h1fd04;
         mem[1498] =  20'h3f644;
         mem[1499] =  20'h58a04;
         mem[1500] =  20'h1dc8a;
         mem[1501] =  20'h0f066;
         mem[1502] =  20'h1dc8a;
         mem[1503] =  20'h1948a;
         mem[1504] =  20'h35c87;
         mem[1505] =  20'h33487;
         mem[1506] =  20'h6cca4;
         mem[1507] =  20'h650e3;
         mem[1508] =  20'h70b05;
         mem[1509] =  20'h0e88b;
         mem[1510] =  20'h10088;
         mem[1511] =  20'h0c983;
         mem[1512] =  20'h14583;
         mem[1513] =  20'h0ccc6;
         mem[1514] =  20'h368c3;
         mem[1515] =  20'h13c85;
         mem[1516] =  20'h8b241;
         mem[1517] =  20'h45241;
         mem[1518] =  20'h452c1;
         mem[1519] =  20'h45583;
         mem[1520] =  20'h368c3;
         mem[1521] =  20'h320c3;
         mem[1522] =  20'h60c49;
         mem[1523] =  20'h5f922;
         mem[1524] =  20'h59ce6;
         mem[1525] =  20'h53066;
         mem[1526] =  20'h60cc4;
         mem[1527] =  20'h1ac50;
         mem[1528] =  20'h60c49;
         mem[1529] =  20'h60449;
         mem[1530] =  20'h488c5;
         mem[1531] =  20'h32dc2;
         mem[1532] =  20'h26a24;
         mem[1533] =  20'h39d87;
         mem[1534] =  20'h1b123;
         mem[1535] =  20'h2ed83;
         mem[1536] =  20'h47925;
         mem[1537] =  20'h4ba41;
         mem[1538] =  20'h72922;
         mem[1539] =  20'h0c922;
         mem[1540] =  20'h51702;
         mem[1541] =  20'h4ba83;
         mem[1542] =  20'h22506;
         mem[1543] =  20'h2e485;
         mem[1544] =  20'h21142;
         mem[1545] =  20'h790c4;
         mem[1546] =  20'h238e5;
         mem[1547] =  20'h1f4e5;
         mem[1548] =  20'h0b066;
         mem[1549] =  20'h19664;
         mem[1550] =  20'h1c122;
         mem[1551] =  20'h19d22;
         mem[1552] =  20'h1c142;
         mem[1553] =  20'h1c122;
         mem[1554] =  20'h09449;
         mem[1555] =  20'h08c49;
         mem[1556] =  20'h22c85;
         mem[1557] =  20'h1b88d;
         mem[1558] =  20'h22866;
         mem[1559] =  20'h210c3;
         mem[1560] =  20'h2d942;
         mem[1561] =  20'h024e5;
         mem[1562] =  20'h44d23;
         mem[1563] =  20'h28449;
         mem[1564] =  20'h13867;
         mem[1565] =  20'h744c3;
         mem[1566] =  20'h32943;
         mem[1567] =  20'h1c542;
         mem[1568] =  20'h45ca6;
         mem[1569] =  20'h1e049;
         mem[1570] =  20'h53507;
         mem[1571] =  20'h09583;
         mem[1572] =  20'h19849;
         mem[1573] =  20'h2ca41;
         mem[1574] =  20'h77a02;
         mem[1575] =  20'h3b8c3;
         mem[1576] =  20'h26ce3;
         mem[1577] =  20'h23885;
         mem[1578] =  20'h13681;
         mem[1579] =  20'h0f866;
         mem[1580] =  20'h28049;
         mem[1581] =  20'h15c4b;
         mem[1582] =  20'h1544b;
         mem[1583] =  20'h15c85;
         mem[1584] =  20'h09432;
         mem[1585] =  20'h0f866;
         mem[1586] =  20'h12e61;
         mem[1587] =  20'h66522;
         mem[1588] =  20'h33cc5;
         mem[1589] =  20'h03849;
         mem[1590] =  20'h02049;
         mem[1591] =  20'h48085;
         mem[1592] =  20'h25e41;
         mem[1593] =  20'h3a9c2;
         mem[1594] =  20'h6ae41;
         mem[1595] =  20'h7a922;
         mem[1596] =  20'h320c3;
         mem[1597] =  20'h6c8e4;
         mem[1598] =  20'h71281;
         mem[1599] =  20'h7a922;
         mem[1600] =  20'h0d9e2;
         mem[1601] =  20'h238c3;
         mem[1602] =  20'h258c3;
         mem[1603] =  20'h7a922;
         mem[1604] =  20'h76d22;
         mem[1605] =  20'h744c3;
         mem[1606] =  20'h714c3;
         mem[1607] =  20'h56485;
         mem[1608] =  20'h59904;
         mem[1609] =  20'h73c66;
         mem[1610] =  20'h51485;
         mem[1611] =  20'h6a703;
         mem[1612] =  20'h0dcc4;
         mem[1613] =  20'h3b066;
         mem[1614] =  20'h20602;
         mem[1615] =  20'h2e485;
         mem[1616] =  20'h340a4;
         mem[1617] =  20'h3b124;
         mem[1618] =  20'h39524;
         mem[1619] =  20'h3bcc3;
         mem[1620] =  20'h32a84;
         mem[1621] =  20'h4c228;
         mem[1622] =  20'h408e3;
         mem[1623] =  20'h3eee1;
         mem[1624] =  20'h02449;
         mem[1625] =  20'h16049;
         mem[1626] =  20'h08c4d;
         mem[1627] =  20'h90e41;
         mem[1628] =  20'h40066;
         mem[1629] =  20'h03838;
         mem[1630] =  20'h02438;
         mem[1631] =  20'h0ecca;
         mem[1632] =  20'h538a6;
         mem[1633] =  20'h858c3;
         mem[1634] =  20'h0904b;
         mem[1635] =  20'h2e0a4;
         mem[1636] =  20'h030b2;
         mem[1637] =  20'h09c50;
         mem[1638] =  20'h08450;
         mem[1639] =  20'h23cc3;
         mem[1640] =  20'h26641;
         mem[1641] =  20'h23cc3;
         mem[1642] =  20'h1f4c3;
         mem[1643] =  20'h54962;
         mem[1644] =  20'h2e4a4;
         mem[1645] =  20'h3b0a7;
         mem[1646] =  20'h3a4a7;
         mem[1647] =  20'h1d066;
         mem[1648] =  20'h26ca4;
         mem[1649] =  20'h85103;
         mem[1650] =  20'h85903;
         mem[1651] =  20'h22967;
         mem[1652] =  20'h3f485;
         mem[1653] =  20'h05066;
         mem[1654] =  20'h0e452;
         mem[1655] =  20'h03c49;
         mem[1656] =  20'h5dce3;
         mem[1657] =  20'h56085;
         mem[1658] =  20'h00466;
         mem[1659] =  20'h2ec66;
         mem[1660] =  20'h51885;
         mem[1661] =  20'h8a661;
         mem[1662] =  20'h14c4d;
         mem[1663] =  20'h46241;
         mem[1664] =  20'h2e0a4;
         mem[1665] =  20'h2e885;
         mem[1666] =  20'h13e02;
         mem[1667] =  20'h07e41;
         mem[1668] =  20'h078a4;
         mem[1669] =  20'h74cc3;
         mem[1670] =  20'h608c3;
         mem[1671] =  20'h3ed64;
         mem[1672] =  20'h3ac66;
         mem[1673] =  20'h47485;
         mem[1674] =  20'h2e8a7;
         mem[1675] =  20'h0f48a;
         mem[1676] =  20'h0ec8a;
         mem[1677] =  20'h1cd23;
         mem[1678] =  20'h32143;
         mem[1679] =  20'h38ea2;
         mem[1680] =  20'h19168;
         mem[1681] =  20'h470cb;
         mem[1682] =  20'h2e066;
         mem[1683] =  20'h048c9;
         mem[1684] =  20'h000c9;
         mem[1685] =  20'h09562;
         mem[1686] =  20'h0d642;
         mem[1687] =  20'h2c6c2;
         mem[1688] =  20'h140c3;
         mem[1689] =  20'h5a849;
         mem[1690] =  20'h5a049;
         mem[1691] =  20'h78241;
         mem[1692] =  20'h0246d;
         mem[1693] =  20'h1acc4;
         mem[1694] =  20'h0ec86;
         mem[1695] =  20'h0da41;
         mem[1696] =  20'h4b0c4;
         mem[1697] =  20'h60849;
         mem[1698] =  20'h4144d;
         mem[1699] =  20'h72241;
         mem[1700] =  20'h1bc49;
         mem[1701] =  20'h03049;
         mem[1702] =  20'h26ca4;
         mem[1703] =  20'h54ca4;
         mem[1704] =  20'h528a4;
         mem[1705] =  20'h54d22;
         mem[1706] =  20'h2bee5;
         mem[1707] =  20'h29906;
         mem[1708] =  20'h718c3;
         mem[1709] =  20'h7f122;
         mem[1710] =  20'h70a41;
         mem[1711] =  20'h54962;
         mem[1712] =  20'h51562;
         mem[1713] =  20'h3b583;
         mem[1714] =  20'h7e904;
         mem[1715] =  20'h731c2;
         mem[1716] =  20'h0cea1;
         mem[1717] =  20'h0c983;
         mem[1718] =  20'h5f485;
         mem[1719] =  20'h470e3;
         mem[1720] =  20'h70cc3;
         mem[1721] =  20'h79485;
         mem[1722] =  20'h4cc85;
         mem[1723] =  20'h4d4c4;
         mem[1724] =  20'h08c66;
         mem[1725] =  20'h5ea61;
         mem[1726] =  20'h2d8a5;
         mem[1727] =  20'h4bd2c;
         mem[1728] =  20'h0284c;
         mem[1729] =  20'h13a23;
         mem[1730] =  20'h0288b;
         mem[1731] =  20'h0106d;
         mem[1732] =  20'h46203;
         mem[1733] =  20'h598a6;
         mem[1734] =  20'h858c3;
         mem[1735] =  20'h00c66;
         mem[1736] =  20'h06e81;
         mem[1737] =  20'h27caa;
         mem[1738] =  20'h28449;
         mem[1739] =  20'h02c49;
         mem[1740] =  20'h04049;
         mem[1741] =  20'h72522;
         mem[1742] =  20'h04049;
         mem[1743] =  20'h01849;
         mem[1744] =  20'h0b050;
         mem[1745] =  20'h07050;
         mem[1746] =  20'h678c3;
         mem[1747] =  20'h12cc3;
         mem[1748] =  20'h21866;
         mem[1749] =  20'h40066;
         mem[1750] =  20'h61468;
         mem[1751] =  20'h3f8e6;
         mem[1752] =  20'h33d82;
         mem[1753] =  20'h0ec54;
         mem[1754] =  20'h678c3;
         mem[1755] =  20'h28849;
         mem[1756] =  20'h678c3;
         mem[1757] =  20'h8adc2;
         mem[1758] =  20'h3fa06;
         mem[1759] =  20'h28449;
         mem[1760] =  20'h0d6a2;
         mem[1761] =  20'h650c3;
         mem[1762] =  20'h810a4;
         mem[1763] =  20'h01108;
         mem[1764] =  20'h28ce3;
         mem[1765] =  20'h41085;
         mem[1766] =  20'h618c4;
         mem[1767] =  20'h2ecc4;
         mem[1768] =  20'h288e3;
         mem[1769] =  20'h26525;
         mem[1770] =  20'h030d5;
         mem[1771] =  20'h02115;
         mem[1772] =  20'h78641;
         mem[1773] =  20'h6a522;
         mem[1774] =  20'h1a261;
         mem[1775] =  20'h19301;
         mem[1776] =  20'h67d22;
         mem[1777] =  20'h64122;
         mem[1778] =  20'h65a41;
         mem[1779] =  20'h71641;
         mem[1780] =  20'h03437;
         mem[1781] =  20'h14503;
         mem[1782] =  20'h6be41;
         mem[1783] =  20'h02837;
         mem[1784] =  20'h4d885;
         mem[1785] =  20'h4cd44;
         mem[1786] =  20'h3c867;
         mem[1787] =  20'h13543;
         mem[1788] =  20'h2e8a6;
         mem[1789] =  20'h194c5;
         mem[1790] =  20'h16922;
         mem[1791] =  20'h0cc85;
         mem[1792] =  20'h21ca4;
         mem[1793] =  20'h02cf8;
         mem[1794] =  20'h78942;
         mem[1795] =  20'h79485;
         mem[1796] =  20'h61849;
         mem[1797] =  20'h8a641;
         mem[1798] =  20'h61849;
         mem[1799] =  20'h5f849;
         mem[1800] =  20'h28849;
         mem[1801] =  20'h1504b;
         mem[1802] =  20'h16922;
         mem[1803] =  20'h335c4;
         mem[1804] =  20'h1b1e3;
         mem[1805] =  20'h0e485;
         mem[1806] =  20'h0f86c;
         mem[1807] =  20'h0ec6c;
         mem[1808] =  20'h2d8c4;
         mem[1809] =  20'h1548a;
         mem[1810] =  20'h28d03;
         mem[1811] =  20'h088c9;
         mem[1812] =  20'h344c5;
         mem[1813] =  20'h0018b;
         mem[1814] =  20'h74122;
         mem[1815] =  20'h7d304;
         mem[1816] =  20'h79d62;
         mem[1817] =  20'h70d22;
         mem[1818] =  20'h33ca4;
         mem[1819] =  20'h60849;
         mem[1820] =  20'h748c3;
         mem[1821] =  20'h710c3;
         mem[1822] =  20'h27a03;
         mem[1823] =  20'h2bd42;
         mem[1824] =  20'h26e41;
         mem[1825] =  20'h38d23;
         mem[1826] =  20'h22d43;
         mem[1827] =  20'h2ca41;
         mem[1828] =  20'h1b5e2;
         mem[1829] =  20'h3f9e2;
         mem[1830] =  20'h22582;
         mem[1831] =  20'h3444c;
         mem[1832] =  20'h03449;
         mem[1833] =  20'h4b066;
         mem[1834] =  20'h5b142;
         mem[1835] =  20'h3f243;
         mem[1836] =  20'h6d143;
         mem[1837] =  20'h274a4;
         mem[1838] =  20'h28ce3;
         mem[1839] =  20'h53067;
         mem[1840] =  20'h42c66;
         mem[1841] =  20'h3f866;
         mem[1842] =  20'h3b886;
         mem[1843] =  20'h1544e;
         mem[1844] =  20'h04832;
         mem[1845] =  20'h4e10c;
         mem[1846] =  20'h0444e;
         mem[1847] =  20'h0144e;
         mem[1848] =  20'h10894;
         mem[1849] =  20'h0d894;
         mem[1850] =  20'h04851;
         mem[1851] =  20'h01051;
         mem[1852] =  20'h35d22;
         mem[1853] =  20'h32122;
         mem[1854] =  20'h0b44d;
         mem[1855] =  20'h06c4d;
         mem[1856] =  20'h04049;
         mem[1857] =  20'h40c87;
         mem[1858] =  20'h47d82;
         mem[1859] =  20'h44d82;
         mem[1860] =  20'h3fdc3;
         mem[1861] =  20'h64281;
         mem[1862] =  20'h41885;
         mem[1863] =  20'h2d1a3;
         mem[1864] =  20'h348c6;
         mem[1865] =  20'h02049;
         mem[1866] =  20'h46582;
         mem[1867] =  20'h265e4;
         mem[1868] =  20'h04085;
         mem[1869] =  20'h5f4c3;
         mem[1870] =  20'h59905;
         mem[1871] =  20'h07c32;
         mem[1872] =  20'h0284e;
         mem[1873] =  20'h15849;
         mem[1874] =  20'h100c3;
         mem[1875] =  20'h25a22;
         mem[1876] =  20'h810a4;
         mem[1877] =  20'h7dca4;
         mem[1878] =  20'h78641;
         mem[1879] =  20'h01085;
         mem[1880] =  20'h17066;
         mem[1881] =  20'h4b84c;
         mem[1882] =  20'h19aa1;
         mem[1883] =  20'h13c66;
         mem[1884] =  20'h368c3;
         mem[1885] =  20'h5fd09;
         mem[1886] =  20'h52d25;
         mem[1887] =  20'h270a6;
         mem[1888] =  20'h3bc66;
         mem[1889] =  20'h020ab;
         mem[1890] =  20'h3c066;
         mem[1891] =  20'h39c66;
         mem[1892] =  20'h22ca4;
         mem[1893] =  20'h1a104;
         mem[1894] =  20'h2d8c3;
         mem[1895] =  20'h0206d;
         mem[1896] =  20'h03449;
         mem[1897] =  20'h02449;
         mem[1898] =  20'h1b143;
         mem[1899] =  20'h12e41;
         mem[1900] =  20'h558e3;
         mem[1901] =  20'h514e3;
         mem[1902] =  20'h11c35;
         mem[1903] =  20'h514a4;
         mem[1904] =  20'h35182;
         mem[1905] =  20'h38a81;
         mem[1906] =  20'h33661;
         mem[1907] =  20'h57d22;
         mem[1908] =  20'h591c4;
         mem[1909] =  20'h4c5c6;
         mem[1910] =  20'h4e867;
         mem[1911] =  20'h6aa42;
         mem[1912] =  20'h6d0c3;
         mem[1913] =  20'h32122;
         mem[1914] =  20'h41d43;
         mem[1915] =  20'h3ed43;
         mem[1916] =  20'h38582;
         mem[1917] =  20'h4b544;
         mem[1918] =  20'h4e867;
         mem[1919] =  20'h4cc67;
         mem[1920] =  20'h4e085;
         mem[1921] =  20'h4d085;
         mem[1922] =  20'h41c4a;
         mem[1923] =  20'h60942;
         mem[1924] =  20'h40c66;
         mem[1925] =  20'h080e3;
         mem[1926] =  20'h2d5a3;
         mem[1927] =  20'h21c85;
         mem[1928] =  20'h4d942;
         mem[1929] =  20'h658a4;
         mem[1930] =  20'h03c49;
         mem[1931] =  20'h408c6;
         mem[1932] =  20'h1bd22;
         mem[1933] =  20'h7f0e3;
         mem[1934] =  20'h452c1;
         mem[1935] =  20'h70a41;
         mem[1936] =  20'h03c49;
         mem[1937] =  20'h01c49;
         mem[1938] =  20'h11854;
         mem[1939] =  20'h0d054;
         mem[1940] =  20'h2f467;
         mem[1941] =  20'h06c49;
         mem[1942] =  20'h67122;
         mem[1943] =  20'h5e122;
         mem[1944] =  20'h33de2;
         mem[1945] =  20'h34066;
         mem[1946] =  20'h288c3;
         mem[1947] =  20'h77542;
         mem[1948] =  20'h740c3;
         mem[1949] =  20'h20127;
         mem[1950] =  20'h29c49;
         mem[1951] =  20'h26c49;
         mem[1952] =  20'h03449;
         mem[1953] =  20'h02449;
         mem[1954] =  20'h22849;
         mem[1955] =  20'h22466;
         mem[1956] =  20'h09503;
         mem[1957] =  20'h5404b;
         mem[1958] =  20'h0b466;
         mem[1959] =  20'h70e41;
         mem[1960] =  20'h6c144;
         mem[1961] =  20'h7e942;
         mem[1962] =  20'h66522;
         mem[1963] =  20'h06866;
         mem[1964] =  20'h36ca4;
         mem[1965] =  20'h01088;
         mem[1966] =  20'h26661;
         mem[1967] =  20'h1f8c3;
         mem[1968] =  20'h088e8;
         mem[1969] =  20'h20604;
         mem[1970] =  20'h07e41;
         mem[1971] =  20'h45d47;
         mem[1972] =  20'h48885;
         mem[1973] =  20'h72cc3;
         mem[1974] =  20'h73886;
         mem[1975] =  20'h5f469;
         mem[1976] =  20'h488c4;
         mem[1977] =  20'h458c4;
         mem[1978] =  20'h3bd23;
         mem[1979] =  20'h5e182;
         mem[1980] =  20'h6dd42;
         mem[1981] =  20'h6a542;
         mem[1982] =  20'h67cc3;
         mem[1983] =  20'h64cc3;
         mem[1984] =  20'h21888;
         mem[1985] =  20'h70cc3;
         mem[1986] =  20'h86942;
         mem[1987] =  20'h83942;
         mem[1988] =  20'h7ea41;
         mem[1989] =  20'h78c85;
         mem[1990] =  20'h0cb02;
         mem[1991] =  20'h190c3;
         mem[1992] =  20'h3bd43;
         mem[1993] =  20'h77264;
         mem[1994] =  20'h10142;
         mem[1995] =  20'h408ee;
         mem[1996] =  20'h41088;
         mem[1997] =  20'h34ca4;
         mem[1998] =  20'h21c49;
         mem[1999] =  20'h2184a;
         mem[2000] =  20'h1c84d;
         mem[2001] =  20'h1b04d;
         mem[2002] =  20'h2e866;
         mem[2003] =  20'h26503;
         mem[2004] =  20'h1c507;
         mem[2005] =  20'h00182;
         mem[2006] =  20'h09466;
         mem[2007] =  20'h090e4;
         mem[2008] =  20'h6cce3;
         mem[2009] =  20'h14c85;
         mem[2010] =  20'h15885;
         mem[2011] =  20'h0f04d;
         mem[2012] =  20'h0f833;
         mem[2013] =  20'h2e466;
         mem[2014] =  20'h8a942;
         mem[2015] =  20'h64182;
         mem[2016] =  20'h15885;
         mem[2017] =  20'h3ec87;
         mem[2018] =  20'h798c3;
         mem[2019] =  20'h018ac;
         mem[2020] =  20'h22ce7;
         mem[2021] =  20'h33ca4;
         mem[2022] =  20'h09466;
         mem[2023] =  20'h28983;
         mem[2024] =  20'h15885;
         mem[2025] =  20'h51962;
         mem[2026] =  20'h59d82;
         mem[2027] =  20'h2bd22;
         mem[2028] =  20'h2c2e2;
         mem[2029] =  20'h3ee64;
         mem[2030] =  20'h344c7;
         mem[2031] =  20'h790c3;
         mem[2032] =  20'h5a449;
         mem[2033] =  20'h2844c;
         mem[2034] =  20'h04849;
         mem[2035] =  20'h01049;
         mem[2036] =  20'h0a04b;
         mem[2037] =  20'h57d06;
         mem[2038] =  20'h420e3;
         mem[2039] =  20'h4bd22;
         mem[2040] =  20'h0a04b;
         mem[2041] =  20'h0804b;
         mem[2042] =  20'h2f542;
         mem[2043] =  20'h41867;
         mem[2044] =  20'h2d8a4;
         mem[2045] =  20'h32085;
         mem[2046] =  20'h04c86;
         mem[2047] =  20'h00486;
         mem[2048] =  20'h23450;
         mem[2049] =  20'h20c50;
         mem[2050] =  20'h04450;
         mem[2051] =  20'h01450;
         mem[2052] =  20'h12f01;
         mem[2053] =  20'h14942;
         mem[2054] =  20'h196e4;
         mem[2055] =  20'h70e61;
         mem[2056] =  20'h78641;
         mem[2057] =  20'h77122;
         mem[2058] =  20'h744c3;
         mem[2059] =  20'h714c3;
         mem[2060] =  20'h6b683;
         mem[2061] =  20'h3e867;
         mem[2062] =  20'h78641;
         mem[2063] =  20'h4cc67;
         mem[2064] =  20'h418c5;
         mem[2065] =  20'h400c5;
         mem[2066] =  20'h0ecc9;
         mem[2067] =  20'h268a5;
         mem[2068] =  20'h5c849;
         mem[2069] =  20'h58049;
         mem[2070] =  20'h0984a;
         mem[2071] =  20'h864c3;
         mem[2072] =  20'h0984a;
         mem[2073] =  20'h644a4;
         mem[2074] =  20'h0984a;
         mem[2075] =  20'h00833;
         mem[2076] =  20'h0984a;
         mem[2077] =  20'h06c49;
         mem[2078] =  20'h39262;
         mem[2079] =  20'h65d22;
         mem[2080] =  20'h1d4e3;
         mem[2081] =  20'h1a5c4;
         mem[2082] =  20'h1d103;
         mem[2083] =  20'h19103;
         mem[2084] =  20'h03d22;
         mem[2085] =  20'h64122;
         mem[2086] =  20'h2e0c8;
         mem[2087] =  20'h45c49;
         mem[2088] =  20'h22449;
         mem[2089] =  20'h28049;
         mem[2090] =  20'h0984a;
         mem[2091] =  20'h0884a;
         mem[2092] =  20'h3bd23;
         mem[2093] =  20'h1b049;
         mem[2094] =  20'h66886;
         mem[2095] =  20'h00124;
         mem[2096] =  20'h228e6;
         mem[2097] =  20'h150a7;
         mem[2098] =  20'h5b142;
         mem[2099] =  20'h64085;
         mem[2100] =  20'h452c1;
         mem[2101] =  20'h3ac4a;
         mem[2102] =  20'h10866;
         mem[2103] =  20'h28049;
         mem[2104] =  20'h350a8;
         mem[2105] =  20'h08486;
         mem[2106] =  20'h098c7;
         mem[2107] =  20'h64982;
         mem[2108] =  20'h798c3;
         mem[2109] =  20'h788c3;
         mem[2110] =  20'h1c44a;
         mem[2111] =  20'h7d261;
         mem[2112] =  20'h4e0c4;
         mem[2113] =  20'h4d10b;
         mem[2114] =  20'h4e0c4;
         mem[2115] =  20'h4c8c4;
         mem[2116] =  20'h358c3;
         mem[2117] =  20'h32302;
         mem[2118] =  20'h5b142;
         mem[2119] =  20'h57942;
         mem[2120] =  20'h2ce61;
         mem[2121] =  20'h2c261;
         mem[2122] =  20'h13e03;
         mem[2123] =  20'h08505;
         mem[2124] =  20'h458c5;
         mem[2125] =  20'h28449;
         mem[2126] =  20'h70a41;
         mem[2127] =  20'h91641;
         mem[2128] =  20'h5e4c3;
         mem[2129] =  20'h624c3;
         mem[2130] =  20'h5dcc3;
         mem[2131] =  20'h79885;
         mem[2132] =  20'h59cc8;
         mem[2133] =  20'h4cd45;
         mem[2134] =  20'h1384d;
         mem[2135] =  20'h0ac6d;
         mem[2136] =  20'h08049;
         mem[2137] =  20'h1106b;
         mem[2138] =  20'h0d46b;
         mem[2139] =  20'h59de2;
         mem[2140] =  20'h13681;
         mem[2141] =  20'h28049;
         mem[2142] =  20'h26cc7;
         mem[2143] =  20'h02c49;
         mem[2144] =  20'h02866;
         mem[2145] =  20'h28849;
         mem[2146] =  20'h074ca;
         mem[2147] =  20'h2d523;
         mem[2148] =  20'h2e123;
         mem[2149] =  20'h7f4c3;
         mem[2150] =  20'h28449;
         mem[2151] =  20'h0f08f;
         mem[2152] =  20'h19a41;
         mem[2153] =  20'h1e449;
         mem[2154] =  20'h0ca61;
         mem[2155] =  20'h0dde2;
         mem[2156] =  20'h0f8e5;
         mem[2157] =  20'h0cd6e;
         mem[2158] =  20'h60449;
         mem[2159] =  20'h72241;
         mem[2160] =  20'h4d466;
         mem[2161] =  20'h06e81;
         mem[2162] =  20'h334a4;
         mem[2163] =  20'h28885;
         mem[2164] =  20'h4d466;
         mem[2165] =  20'h5c085;
         mem[2166] =  20'h58085;
         mem[2167] =  20'h748c3;
         mem[2168] =  20'h25cc3;
         mem[2169] =  20'h15c34;
         mem[2170] =  20'h268e3;
         mem[2171] =  20'h21c8d;
         mem[2172] =  20'h39885;
         mem[2173] =  20'h678a4;
         mem[2174] =  20'h33c67;
         mem[2175] =  20'h33d42;
         mem[2176] =  20'h26241;
         mem[2177] =  20'h209e4;
         mem[2178] =  20'h40509;
         mem[2179] =  20'h44f01;
         mem[2180] =  20'h0d04d;
         mem[2181] =  20'h05085;
         mem[2182] =  20'h1a543;
         mem[2183] =  20'h2d241;
         mem[2184] =  20'h0cb01;
         mem[2185] =  20'h1c44b;
         mem[2186] =  20'h00085;
         mem[2187] =  20'h6b641;
         mem[2188] =  20'h6ae41;
         mem[2189] =  20'h03125;
         mem[2190] =  20'h15d55;
         mem[2191] =  20'h2d4e3;
         mem[2192] =  20'h384c3;
         mem[2193] =  20'h5a0e4;
         mem[2194] =  20'h594e4;
         mem[2195] =  20'h860c3;
         mem[2196] =  20'h850c3;
         mem[2197] =  20'h1e449;
         mem[2198] =  20'h32e41;
         mem[2199] =  20'h1e449;
         mem[2200] =  20'h6c142;
         mem[2201] =  20'h66563;
         mem[2202] =  20'h44c85;
         mem[2203] =  20'h74522;
         mem[2204] =  20'h1f849;
         mem[2205] =  20'h35485;
         mem[2206] =  20'h33c85;
         mem[2207] =  20'h35485;
         mem[2208] =  20'h34867;
         mem[2209] =  20'h35485;
         mem[2210] =  20'h28067;
         mem[2211] =  20'h35485;
         mem[2212] =  20'h47486;
         mem[2213] =  20'h461c6;
         mem[2214] =  20'h12d62;
         mem[2215] =  20'h4144a;
         mem[2216] =  20'h77562;
         mem[2217] =  20'h74522;
         mem[2218] =  20'h45241;
         mem[2219] =  20'h1b88d;
         mem[2220] =  20'h76e41;
         mem[2221] =  20'h78641;
         mem[2222] =  20'h70922;
         mem[2223] =  20'h6d922;
         mem[2224] =  20'h6ad22;
         mem[2225] =  20'h09870;
         mem[2226] =  20'h08470;
         mem[2227] =  20'h2284a;
         mem[2228] =  20'h2184a;
         mem[2229] =  20'h03058;
         mem[2230] =  20'h19c4a;
         mem[2231] =  20'h04049;
         mem[2232] =  20'h01849;
         mem[2233] =  20'h21cc5;
         mem[2234] =  20'h27449;
         mem[2235] =  20'h0f8a8;
         mem[2236] =  20'h0e4a8;
         mem[2237] =  20'h02849;
         mem[2238] =  20'h19c66;
         mem[2239] =  20'h04092;
         mem[2240] =  20'h01092;
         mem[2241] =  20'h38702;
         mem[2242] =  20'h2e8e3;
         mem[2243] =  20'h3488f;
         mem[2244] =  20'h030ae;
         mem[2245] =  20'h42c85;
         mem[2246] =  20'h01449;
         mem[2247] =  20'h0a468;
         mem[2248] =  20'h07868;
         mem[2249] =  20'h3f644;
         mem[2250] =  20'h58a02;
         mem[2251] =  20'h58a05;
         mem[2252] =  20'h3f485;
         mem[2253] =  20'h74903;
         mem[2254] =  20'h65885;
         mem[2255] =  20'h67922;
         mem[2256] =  20'h65d22;
         mem[2257] =  20'h58a04;
         mem[2258] =  20'h5de62;
         mem[2259] =  20'h60522;
         mem[2260] =  20'h01837;
         mem[2261] =  20'h3eb02;
         mem[2262] =  20'h384a4;
         mem[2263] =  20'h39269;
         mem[2264] =  20'h47066;
         mem[2265] =  20'h22584;
         mem[2266] =  20'h7e922;
         mem[2267] =  20'h40942;
         mem[2268] =  20'h32a81;
         mem[2269] =  20'h418ea;
         mem[2270] =  20'h3fcea;
         mem[2271] =  20'h48449;
         mem[2272] =  20'h348ac;
         mem[2273] =  20'h3b4c4;
         mem[2274] =  20'h59467;
         mem[2275] =  20'h10cc8;
         mem[2276] =  20'h02449;
         mem[2277] =  20'h67522;
         mem[2278] =  20'h4b162;
         mem[2279] =  20'h4e163;
         mem[2280] =  20'h27c66;
         mem[2281] =  20'h02849;
         mem[2282] =  20'h344c7;
         mem[2283] =  20'h32302;
         mem[2284] =  20'h46d0a;
         mem[2285] =  20'h150d5;
         mem[2286] =  20'h4d44a;
         mem[2287] =  20'h67ca4;
         mem[2288] =  20'h28049;
         mem[2289] =  20'h42466;
         mem[2290] =  20'h40066;
         mem[2291] =  20'h4fc66;
         mem[2292] =  20'h4b866;
         mem[2293] =  20'h60c49;
         mem[2294] =  20'h60449;
         mem[2295] =  20'h808a4;
         mem[2296] =  20'h7e4a4;
         mem[2297] =  20'h79922;
         mem[2298] =  20'h19dc2;
         mem[2299] =  20'h15542;
         mem[2300] =  20'h5f0a4;
         mem[2301] =  20'h11833;
         mem[2302] =  20'h4cc68;
         mem[2303] =  20'h45ca4;
         mem[2304] =  20'h08503;
         mem[2305] =  20'h40182;
         mem[2306] =  20'h1784a;
         mem[2307] =  20'h26466;
         mem[2308] =  20'h05056;
         mem[2309] =  20'h00856;
         mem[2310] =  20'h65661;
         mem[2311] =  20'h4d885;
         mem[2312] =  20'h28449;
         mem[2313] =  20'h89a41;
         mem[2314] =  20'h33d45;
         mem[2315] =  20'h32641;
         mem[2316] =  20'h0f466;
         mem[2317] =  20'h6a707;
         mem[2318] =  20'h3c885;
         mem[2319] =  20'h22449;
         mem[2320] =  20'h3c885;
         mem[2321] =  20'h468a5;
         mem[2322] =  20'h54922;
         mem[2323] =  20'h06661;
         mem[2324] =  20'h72906;
         mem[2325] =  20'h4c908;
         mem[2326] =  20'h40542;
         mem[2327] =  20'h258c3;
         mem[2328] =  20'h73ce3;
         mem[2329] =  20'h714c3;
         mem[2330] =  20'h6d4c3;
         mem[2331] =  20'h775e4;
         mem[2332] =  20'h59cc8;
         mem[2333] =  20'h400e4;
         mem[2334] =  20'h3bcc3;
         mem[2335] =  20'h6b8c3;
         mem[2336] =  20'h35049;
         mem[2337] =  20'h27049;
         mem[2338] =  20'h3c866;
         mem[2339] =  20'h39466;
         mem[2340] =  20'h6dd22;
         mem[2341] =  20'h7d122;
         mem[2342] =  20'h80522;
         mem[2343] =  20'h7d922;
         mem[2344] =  20'h6be41;
         mem[2345] =  20'h6a641;
         mem[2346] =  20'h11c4b;
         mem[2347] =  20'h0cc4b;
         mem[2348] =  20'h03c38;
         mem[2349] =  20'h7fd04;
         mem[2350] =  20'h28c49;
         mem[2351] =  20'h3a0a7;
         mem[2352] =  20'h3bcc3;
         mem[2353] =  20'h390e3;
         mem[2354] =  20'h1e84a;
         mem[2355] =  20'h3a0c3;
         mem[2356] =  20'h030a7;
         mem[2357] =  20'h09126;
         mem[2358] =  20'h03c38;
         mem[2359] =  20'h02038;
         mem[2360] =  20'h4e467;
         mem[2361] =  20'h4d067;
         mem[2362] =  20'h218d3;
         mem[2363] =  20'h27866;
         mem[2364] =  20'h22466;
         mem[2365] =  20'h64ca4;
         mem[2366] =  20'h560a5;
         mem[2367] =  20'h514a5;
         mem[2368] =  20'h1e84a;
         mem[2369] =  20'h1904a;
         mem[2370] =  20'h2d8a4;
         mem[2371] =  20'h798e4;
         mem[2372] =  20'h474c3;
         mem[2373] =  20'h0cb01;
         mem[2374] =  20'h100ea;
         mem[2375] =  20'h51c49;
         mem[2376] =  20'h03453;
         mem[2377] =  20'h46ce3;
         mem[2378] =  20'h0a10a;
         mem[2379] =  20'h404e9;
         mem[2380] =  20'h798a5;
         mem[2381] =  20'h41466;
         mem[2382] =  20'h0a10a;
         mem[2383] =  20'h0690a;
         mem[2384] =  20'h42866;
         mem[2385] =  20'h3fc66;
         mem[2386] =  20'h288a4;
         mem[2387] =  20'h4c0c3;
         mem[2388] =  20'h2d582;
         mem[2389] =  20'h2e0a5;
         mem[2390] =  20'h10522;
         mem[2391] =  20'h20d65;
         mem[2392] =  20'h54486;
         mem[2393] =  20'h1ad22;
         mem[2394] =  20'h0e1a2;
         mem[2395] =  20'h28049;
         mem[2396] =  20'h35049;
         mem[2397] =  20'h7dd42;
         mem[2398] =  20'h5ee81;
         mem[2399] =  20'h6ad22;
         mem[2400] =  20'h03453;
         mem[2401] =  20'h02453;
         mem[2402] =  20'h1fac1;
         mem[2403] =  20'h0c922;
         mem[2404] =  20'h38709;
         mem[2405] =  20'h26604;
         mem[2406] =  20'h32e42;
         mem[2407] =  20'h0784a;
         mem[2408] =  20'h04066;
         mem[2409] =  20'h01466;
         mem[2410] =  20'h2e485;
         mem[2411] =  20'h20ce5;
         mem[2412] =  20'h0f942;
         mem[2413] =  20'h4ba61;
         mem[2414] =  20'h35049;
         mem[2415] =  20'h34849;
         mem[2416] =  20'h35449;
         mem[2417] =  20'h46469;
         mem[2418] =  20'h3a8c5;
         mem[2419] =  20'h5804a;
         mem[2420] =  20'h80903;
         mem[2421] =  20'h8a641;
         mem[2422] =  20'h1b8a6;
         mem[2423] =  20'h6ad82;
         mem[2424] =  20'h490c3;
         mem[2425] =  20'h4b942;
         mem[2426] =  20'h76f02;
         mem[2427] =  20'h72522;
         mem[2428] =  20'h0a84b;
         mem[2429] =  20'h0784b;
         mem[2430] =  20'h66d03;
         mem[2431] =  20'h08449;
         mem[2432] =  20'h41466;
         mem[2433] =  20'h334c3;
         mem[2434] =  20'h488a4;
         mem[2435] =  20'h45ca4;
         mem[2436] =  20'h29466;
         mem[2437] =  20'h27066;
         mem[2438] =  20'h3b4e4;
         mem[2439] =  20'h34467;
         mem[2440] =  20'h418c4;
         mem[2441] =  20'h20449;
         mem[2442] =  20'h4c206;
         mem[2443] =  20'h58cea;
         mem[2444] =  20'h5b106;
         mem[2445] =  20'h40c67;
         mem[2446] =  20'h22466;
         mem[2447] =  20'h1b832;
         mem[2448] =  20'h1c167;
         mem[2449] =  20'h32a41;
         mem[2450] =  20'h418c4;
         mem[2451] =  20'h21867;
         mem[2452] =  20'h54486;
         mem[2453] =  20'h53486;
         mem[2454] =  20'h5314b;
         mem[2455] =  20'h06834;
         mem[2456] =  20'h54922;
         mem[2457] =  20'h51d22;
         mem[2458] =  20'h6e122;
         mem[2459] =  20'h6a522;
         mem[2460] =  20'h03d2c;
         mem[2461] =  20'h400c4;
         mem[2462] =  20'h3a542;
         mem[2463] =  20'h38923;
         mem[2464] =  20'h2d641;
         mem[2465] =  20'h2e468;
         mem[2466] =  20'h4e04c;
         mem[2467] =  20'h5ea41;
         mem[2468] =  20'h6ec67;
         mem[2469] =  20'h57d42;
         mem[2470] =  20'h6ec67;
         mem[2471] =  20'h15833;
         mem[2472] =  20'h6ec67;
         mem[2473] =  20'h1a963;
         mem[2474] =  20'h6ec67;
         mem[2475] =  20'h33963;
         mem[2476] =  20'h2fc85;
         mem[2477] =  20'h1c153;
         mem[2478] =  20'h088e6;
         mem[2479] =  20'h20cc7;
         mem[2480] =  20'h02c49;
         mem[2481] =  20'h46485;
         mem[2482] =  20'h2fc85;
         mem[2483] =  20'h2cc85;
         mem[2484] =  20'h6ec67;
         mem[2485] =  20'h27885;
         mem[2486] =  20'h62469;
         mem[2487] =  20'h5e869;
         mem[2488] =  20'h42467;
         mem[2489] =  20'h40067;
         mem[2490] =  20'h624a4;
         mem[2491] =  20'h06466;
         mem[2492] =  20'h03466;
         mem[2493] =  20'h01ca6;
         mem[2494] =  20'h07508;
         mem[2495] =  20'h89a61;
         mem[2496] =  20'h3c122;
         mem[2497] =  20'h26522;
         mem[2498] =  20'h27cc5;
         mem[2499] =  20'h3a466;
         mem[2500] =  20'h1a5c3;
         mem[2501] =  20'h00c8a;
         mem[2502] =  20'h140e3;
         mem[2503] =  20'h28085;
         mem[2504] =  20'h0748e;
         mem[2505] =  20'h582c2;
         mem[2506] =  20'h7f0c3;
         mem[2507] =  20'h0ac67;
         mem[2508] =  20'h00c66;
         mem[2509] =  20'h4c226;
         mem[2510] =  20'h018c3;
         mem[2511] =  20'h2f122;
         mem[2512] =  20'h58942;
         mem[2513] =  20'h3b4a6;
         mem[2514] =  20'h08503;
         mem[2515] =  20'h48066;
         mem[2516] =  20'h46c66;
         mem[2517] =  20'h45a61;
         mem[2518] =  20'h1f4c3;
         mem[2519] =  20'h74142;
         mem[2520] =  20'h70942;
         mem[2521] =  20'h61522;
         mem[2522] =  20'h6a641;
         mem[2523] =  20'h6be41;
         mem[2524] =  20'h7d122;
         mem[2525] =  20'h61522;
         mem[2526] =  20'h0e849;
         mem[2527] =  20'h35c4c;
         mem[2528] =  20'h6c504;
         mem[2529] =  20'h7f8c3;
         mem[2530] =  20'h33c4c;
         mem[2531] =  20'h2d8c3;
         mem[2532] =  20'h28849;
         mem[2533] =  20'h7fcc3;
         mem[2534] =  20'h7ecc3;
         mem[2535] =  20'h0b86a;
         mem[2536] =  20'h0646a;
         mem[2537] =  20'h16849;
         mem[2538] =  20'h258c4;
         mem[2539] =  20'h3ccc3;
         mem[2540] =  20'h14849;
         mem[2541] =  20'h04049;
         mem[2542] =  20'h384c3;
         mem[2543] =  20'h1d88a;
         mem[2544] =  20'h1988a;
         mem[2545] =  20'h61522;
         mem[2546] =  20'h5e122;
         mem[2547] =  20'h600c3;
         mem[2548] =  20'h5f122;
         mem[2549] =  20'h07a41;
         mem[2550] =  20'h0f467;
         mem[2551] =  20'h09466;
         mem[2552] =  20'h08866;
         mem[2553] =  20'h288e3;
         mem[2554] =  20'h0f04d;
         mem[2555] =  20'h47cc3;
         mem[2556] =  20'h088cf;
         mem[2557] =  20'h03467;
         mem[2558] =  20'h26603;
         mem[2559] =  20'h2ec66;
         mem[2560] =  20'h2e049;
         mem[2561] =  20'h03458;
         mem[2562] =  20'h02458;
         mem[2563] =  20'h540a4;
         mem[2564] =  20'h6c122;
         mem[2565] =  20'h39a42;
         mem[2566] =  20'h534a4;
         mem[2567] =  20'h77e22;
         mem[2568] =  20'h12d27;
         mem[2569] =  20'h0cb01;
         mem[2570] =  20'h64241;
         mem[2571] =  20'h02c49;
         mem[2572] =  20'h391c6;
         mem[2573] =  20'h2ec66;
         mem[2574] =  20'h02849;
         mem[2575] =  20'h2884a;
         mem[2576] =  20'h01c49;
         mem[2577] =  20'h024e7;
         mem[2578] =  20'h47485;
         mem[2579] =  20'h2e868;
         mem[2580] =  20'h27c69;
         mem[2581] =  20'h5c485;
         mem[2582] =  20'h57c85;
         mem[2583] =  20'h03c85;
         mem[2584] =  20'h01485;
         mem[2585] =  20'h07cc5;
         mem[2586] =  20'h4d922;
         mem[2587] =  20'h35143;
         mem[2588] =  20'h28067;
         mem[2589] =  20'h22c88;
         mem[2590] =  20'h39104;
         mem[2591] =  20'h33ca4;
         mem[2592] =  20'h4cca4;
         mem[2593] =  20'h7a4a4;
         mem[2594] =  20'h01cc9;
         mem[2595] =  20'h1d8a4;
         mem[2596] =  20'h664c4;
         mem[2597] =  20'h2f0a6;
         mem[2598] =  20'h2d4a6;
         mem[2599] =  20'h280c7;
         mem[2600] =  20'h70a41;
         mem[2601] =  20'h71641;
         mem[2602] =  20'h1a04a;
         mem[2603] =  20'h04098;
         mem[2604] =  20'h0208f;
         mem[2605] =  20'h04098;
         mem[2606] =  20'h1acc9;
         mem[2607] =  20'h5b522;
         mem[2608] =  20'h39123;
         mem[2609] =  20'h368c3;
         mem[2610] =  20'h320c3;
         mem[2611] =  20'h2f122;
         mem[2612] =  20'h06cca;
         mem[2613] =  20'h04477;
         mem[2614] =  20'h5e049;
         mem[2615] =  20'h40942;
         mem[2616] =  20'h25943;
         mem[2617] =  20'h4ec85;
         mem[2618] =  20'h19433;
         mem[2619] =  20'h0b432;
         mem[2620] =  20'h07032;
         mem[2621] =  20'h40cc3;
         mem[2622] =  20'h1b4a9;
         mem[2623] =  20'h530e7;
         mem[2624] =  20'h53ce7;
         mem[2625] =  20'h60866;
         mem[2626] =  20'h58885;
         mem[2627] =  20'h79485;
         mem[2628] =  20'h64ca8;
         mem[2629] =  20'h4ed22;
         mem[2630] =  20'h4b122;
         mem[2631] =  20'h40183;
         mem[2632] =  20'h59ca4;
         mem[2633] =  20'h2ec66;
         mem[2634] =  20'h60449;
         mem[2635] =  20'h3c4e3;
         mem[2636] =  20'h08c56;
         mem[2637] =  20'h270e3;
         mem[2638] =  20'h76e61;
         mem[2639] =  20'h04478;
         mem[2640] =  20'h528a6;
         mem[2641] =  20'h290a7;
         mem[2642] =  20'h25c85;
         mem[2643] =  20'h274c5;
         mem[2644] =  20'h2e466;
         mem[2645] =  20'h358e7;
         mem[2646] =  20'h32ce7;
         mem[2647] =  20'h40da2;
         mem[2648] =  20'h0d466;
         mem[2649] =  20'h52e23;
         mem[2650] =  20'h51a23;
         mem[2651] =  20'h42903;
         mem[2652] =  20'h3e903;
         mem[2653] =  20'h3b585;
         mem[2654] =  20'h0e8a8;
         mem[2655] =  20'h0f0c8;
         mem[2656] =  20'h06522;
         mem[2657] =  20'h11c32;
         mem[2658] =  20'h13433;
         mem[2659] =  20'h37050;
         mem[2660] =  20'h32850;
         mem[2661] =  20'h7f162;
         mem[2662] =  20'h27885;
         mem[2663] =  20'h28485;
         mem[2664] =  20'h15066;
         mem[2665] =  20'h274c5;
         mem[2666] =  20'h35067;
         mem[2667] =  20'h0f466;
         mem[2668] =  20'h6c4c3;
         mem[2669] =  20'h0f466;
         mem[2670] =  20'h13d0a;
         mem[2671] =  20'h288a6;
         mem[2672] =  20'h258e4;
         mem[2673] =  20'h79d62;
         mem[2674] =  20'h2ccc4;
         mem[2675] =  20'h47c85;
         mem[2676] =  20'h09049;
         mem[2677] =  20'h03c36;
         mem[2678] =  20'h02036;
         mem[2679] =  20'h2f122;
         mem[2680] =  20'h2e485;
         mem[2681] =  20'h2ec66;
         mem[2682] =  20'h0252d;
         mem[2683] =  20'h04438;
         mem[2684] =  20'h01838;
         mem[2685] =  20'h794a4;
         mem[2686] =  20'h77641;
         mem[2687] =  20'h38e81;
         mem[2688] =  20'h33d22;
         mem[2689] =  20'h2ca65;
         mem[2690] =  20'h32a61;
         mem[2691] =  20'h35d22;
         mem[2692] =  20'h0e8c8;
         mem[2693] =  20'h3ace4;
         mem[2694] =  20'h1ac70;
         mem[2695] =  20'h36870;
         mem[2696] =  20'h32c70;
         mem[2697] =  20'h0504e;
         mem[2698] =  20'h0084e;
         mem[2699] =  20'h04456;
         mem[2700] =  20'h01456;
         mem[2701] =  20'h10894;
         mem[2702] =  20'h0d894;
         mem[2703] =  20'h28449;
         mem[2704] =  20'h03070;
         mem[2705] =  20'h2ec66;
         mem[2706] =  20'h19d23;
         mem[2707] =  20'h22904;
         mem[2708] =  20'h5dd42;
         mem[2709] =  20'h66122;
         mem[2710] =  20'h0ec66;
         mem[2711] =  20'h0b0a4;
         mem[2712] =  20'h2e066;
         mem[2713] =  20'h2d583;
         mem[2714] =  20'h21c86;
         mem[2715] =  20'h07885;
         mem[2716] =  20'h670c4;
         mem[2717] =  20'h58582;
         mem[2718] =  20'h744c3;
         mem[2719] =  20'h650c3;
         mem[2720] =  20'h4dce9;
         mem[2721] =  20'h3a8c3;
         mem[2722] =  20'h1a661;
         mem[2723] =  20'h0d8c3;
         mem[2724] =  20'h28449;
         mem[2725] =  20'h28049;
         mem[2726] =  20'h5b8a5;
         mem[2727] =  20'h584a5;
         mem[2728] =  20'h28ce3;
         mem[2729] =  20'h53467;
         mem[2730] =  20'h66105;
         mem[2731] =  20'h7f943;
         mem[2732] =  20'h46241;
         mem[2733] =  20'h2604a;
         mem[2734] =  20'h0d281;
         mem[2735] =  20'h5404b;
         mem[2736] =  20'h790c4;
         mem[2737] =  20'h600c3;
         mem[2738] =  20'h4c641;
         mem[2739] =  20'h329e2;
         mem[2740] =  20'h07e41;
         mem[2741] =  20'h01832;
         mem[2742] =  20'h17c4a;
         mem[2743] =  20'h1344a;
         mem[2744] =  20'h21c89;
         mem[2745] =  20'h21c89;
         mem[2746] =  20'h13a81;
         mem[2747] =  20'h1a5a2;
         mem[2748] =  20'h300e7;
         mem[2749] =  20'h2bce7;
         mem[2750] =  20'h470a6;
         mem[2751] =  20'h474a6;
         mem[2752] =  20'h4dc66;
         mem[2753] =  20'h6a641;
         mem[2754] =  20'h6be41;
         mem[2755] =  20'h45d25;
         mem[2756] =  20'h3a9e2;
         mem[2757] =  20'h26cc3;
         mem[2758] =  20'h1a983;
         mem[2759] =  20'h3a066;
         mem[2760] =  20'h2e9a2;
         mem[2761] =  20'h47d6d;
         mem[2762] =  20'h494c3;
         mem[2763] =  20'h44cc3;
         mem[2764] =  20'h2bf01;
         mem[2765] =  20'h2bd42;
         mem[2766] =  20'h33a41;
         mem[2767] =  20'h0c942;
         mem[2768] =  20'h05033;
         mem[2769] =  20'h268c8;
         mem[2770] =  20'h2ac49;
         mem[2771] =  20'h25c49;
         mem[2772] =  20'h8a641;
         mem[2773] =  20'h83522;
         mem[2774] =  20'h750c3;
         mem[2775] =  20'h7ed22;
         mem[2776] =  20'h684a4;
         mem[2777] =  20'h648a4;
         mem[2778] =  20'h04ca6;
         mem[2779] =  20'h000a6;
         mem[2780] =  20'h67d22;
         mem[2781] =  20'h64122;
         mem[2782] =  20'h67942;
         mem[2783] =  20'h64142;
         mem[2784] =  20'h78241;
         mem[2785] =  20'h76e41;
         mem[2786] =  20'h22526;
         mem[2787] =  20'h26ce3;
         mem[2788] =  20'h20665;
         mem[2789] =  20'h0d602;
         mem[2790] =  20'h4c10c;
         mem[2791] =  20'h154cf;
         mem[2792] =  20'h1d033;
         mem[2793] =  20'h1ac33;
         mem[2794] =  20'h5bc85;
         mem[2795] =  20'h58485;
         mem[2796] =  20'h4e066;
         mem[2797] =  20'h460c3;
         mem[2798] =  20'h22c85;
         mem[2799] =  20'h1a8c5;
         mem[2800] =  20'h35d25;
         mem[2801] =  20'h32125;
         mem[2802] =  20'h4e066;
         mem[2803] =  20'h5de41;
         mem[2804] =  20'h4e066;
         mem[2805] =  20'h4d466;
         mem[2806] =  20'h5f641;
         mem[2807] =  20'h25a41;
         mem[2808] =  20'h262c1;
         mem[2809] =  20'h01cea;
         mem[2810] =  20'h15cd1;
         mem[2811] =  20'h144d1;
         mem[2812] =  20'h4d10b;
         mem[2813] =  20'h52603;
         mem[2814] =  20'h4e0c4;
         mem[2815] =  20'h5a087;
         mem[2816] =  20'h43067;
         mem[2817] =  20'h3f467;
         mem[2818] =  20'h52e41;
         mem[2819] =  20'h3fd42;
         mem[2820] =  20'h54522;
         mem[2821] =  20'h51522;
         mem[2822] =  20'h0f832;
         mem[2823] =  20'h0f432;
         mem[2824] =  20'h4dc4a;
         mem[2825] =  20'h518c3;
         mem[2826] =  20'h3bd03;
         mem[2827] =  20'h3ed22;
         mem[2828] =  20'h3a202;
         mem[2829] =  20'h06641;
         mem[2830] =  20'h03049;
         mem[2831] =  20'h22466;
         mem[2832] =  20'h28849;
         mem[2833] =  20'h02849;
         mem[2834] =  20'h1b4c3;
         mem[2835] =  20'h13243;
         mem[2836] =  20'h19301;
         mem[2837] =  20'h65922;
         mem[2838] =  20'h3b485;
         mem[2839] =  20'h209a3;
         mem[2840] =  20'h2ce03;
         mem[2841] =  20'h2cdc3;
         mem[2842] =  20'h2dd22;
         mem[2843] =  20'h38a02;
         mem[2844] =  20'h349a3;
         mem[2845] =  20'h325a3;
         mem[2846] =  20'h1c183;
         mem[2847] =  20'h6a943;
         mem[2848] =  20'h71e41;
         mem[2849] =  20'h6a641;
         mem[2850] =  20'h79122;
         mem[2851] =  20'h7d562;
         mem[2852] =  20'h6c503;
         mem[2853] =  20'h46d05;
         mem[2854] =  20'h20a41;
         mem[2855] =  20'h344a5;
         mem[2856] =  20'h338c3;
         mem[2857] =  20'h26123;
         mem[2858] =  20'h28849;
         mem[2859] =  20'h21c66;
         mem[2860] =  20'h5b049;
         mem[2861] =  20'h59849;
         mem[2862] =  20'h0eca6;
         mem[2863] =  20'h0952c;
         mem[2864] =  20'h52a2b;
         mem[2865] =  20'h0d982;
         mem[2866] =  20'h3bd03;
         mem[2867] =  20'h3a8a9;
         mem[2868] =  20'h03849;
         mem[2869] =  20'h02049;
         mem[2870] =  20'h0904c;
         mem[2871] =  20'h461a2;
         mem[2872] =  20'h39a61;
         mem[2873] =  20'h538c4;
         mem[2874] =  20'h5a485;
         mem[2875] =  20'h00867;
         mem[2876] =  20'h0ac67;
         mem[2877] =  20'h07067;
         mem[2878] =  20'h80122;
         mem[2879] =  20'h0144a;
         mem[2880] =  20'h37086;
         mem[2881] =  20'h32086;
         mem[2882] =  20'h55ca4;
         mem[2883] =  20'h518a4;
         mem[2884] =  20'h55085;
         mem[2885] =  20'h52885;
         mem[2886] =  20'h5f604;
         mem[2887] =  20'h5e604;
         mem[2888] =  20'h614e3;
         mem[2889] =  20'h34867;
         mem[2890] =  20'h54922;
         mem[2891] =  20'h52223;
         mem[2892] =  20'h54905;
         mem[2893] =  20'h52105;
         mem[2894] =  20'h5b8a4;
         mem[2895] =  20'h70963;
         mem[2896] =  20'h64184;
         mem[2897] =  20'h800c3;
         mem[2898] =  20'h50466;
         mem[2899] =  20'h4b066;
         mem[2900] =  20'h7a922;
         mem[2901] =  20'h25d65;
         mem[2902] =  20'h7a922;
         mem[2903] =  20'h76e41;
         mem[2904] =  20'h64e61;
         mem[2905] =  20'h57a41;
         mem[2906] =  20'h7a922;
         mem[2907] =  20'h76d22;
         mem[2908] =  20'h79d22;
         mem[2909] =  20'h77922;
         mem[2910] =  20'h10c34;
         mem[2911] =  20'h6a704;
         mem[2912] =  20'h0946b;
     end

endmodule: rect1_rom
