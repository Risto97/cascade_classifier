module featureThreshold_rom
  #(
     parameter W_DATA = 12,
     parameter W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               8'b00000000: data1 <= -12'h081;
               8'b00000001: data1 <=  12'h032;
               8'b00000010: data1 <=  12'h059;
               8'b00000011: data1 <=  12'h017;
               8'b00000100: data1 <=  12'h03d;
               8'b00000101: data1 <=  12'h197;
               8'b00000110: data1 <=  12'h00b;
               8'b00000111: data1 <= -12'h04d;
               8'b00001000: data1 <=  12'h018;
               8'b00001001: data1 <= -12'h056;
               8'b00001010: data1 <=  12'h053;
               8'b00001011: data1 <=  12'h057;
               8'b00001100: data1 <=  12'h177;
               8'b00001101: data1 <=  12'h094;
               8'b00001110: data1 <= -12'h04e;
               8'b00001111: data1 <=  12'h021;
               8'b00010000: data1 <=  12'h04b;
               8'b00010001: data1 <= -12'h01c;
               8'b00010010: data1 <= -12'h028;
               8'b00010011: data1 <=  12'h040;
               8'b00010100: data1 <= -12'h054;
               8'b00010101: data1 <= -12'h233;
               8'b00010110: data1 <=  12'h03a;
               8'b00010111: data1 <=  12'h029;
               8'b00011000: data1 <=  12'h176;
               8'b00011001: data1 <=  12'h11d;
               8'b00011010: data1 <=  12'h081;
               8'b00011011: data1 <=  12'h03a;
               8'b00011100: data1 <=  12'h03b;
               8'b00011101: data1 <= -12'h00c;
               8'b00011110: data1 <=  12'h086;
               8'b00011111: data1 <= -12'h01d;
               8'b00100000: data1 <=  12'h0ce;
               8'b00100001: data1 <=  12'h0c0;
               8'b00100010: data1 <= -12'h11c;
               8'b00100011: data1 <= -12'h0c8;
               8'b00100100: data1 <=  12'h15b;
               8'b00100101: data1 <= -12'h007;
               8'b00100110: data1 <=  12'h1d9;
               8'b00100111: data1 <= -12'h0d2;
               8'b00101000: data1 <= -12'h0ae;
               8'b00101001: data1 <=  12'h5f2;
               8'b00101010: data1 <=  12'h04f;
               8'b00101011: data1 <=  12'h047;
               8'b00101100: data1 <=  12'h0a2;
               8'b00101101: data1 <= -12'h025;
               8'b00101110: data1 <=  12'h007;
               8'b00101111: data1 <=  12'h07b;
               8'b00110000: data1 <= -12'h142;
               8'b00110001: data1 <=  12'h008;
               8'b00110010: data1 <=  12'h06e;
               8'b00110011: data1 <= -12'h0b8;
               8'b00110100: data1 <= -12'h10d;
               8'b00110101: data1 <=  12'h040;
               8'b00110110: data1 <=  12'h254;
               8'b00110111: data1 <=  12'h019;
               8'b00111000: data1 <=  12'h01b;
               8'b00111001: data1 <=  12'h04b;
               8'b00111010: data1 <=  12'h051;
               8'b00111011: data1 <= -12'h470;
               8'b00111100: data1 <=  12'h025;
               8'b00111101: data1 <= -12'h09a;
               8'b00111110: data1 <=  12'h04b;
               8'b00111111: data1 <= -12'h02d;
               8'b01000000: data1 <=  12'h08a;
               8'b01000001: data1 <= -12'h092;
               8'b01000010: data1 <= -12'h02e;
               8'b01000011: data1 <= -12'h10b;
               8'b01000100: data1 <= -12'h0ad;
               8'b01000101: data1 <=  12'h007;
               8'b01000110: data1 <= -12'h211;
               8'b01000111: data1 <=  12'h05d;
               8'b01001000: data1 <= -12'h08b;
               8'b01001001: data1 <=  12'h06b;
               8'b01001010: data1 <=  12'h05b;
               8'b01001011: data1 <= -12'h017;
               8'b01001100: data1 <=  12'h0b2;
               8'b01001101: data1 <=  12'h0ea;
               8'b01001110: data1 <=  12'h009;
               8'b01001111: data1 <=  12'h035;
               8'b01010000: data1 <= -12'h06c;
               8'b01010001: data1 <= -12'h017;
               8'b01010010: data1 <= -12'h043;
               8'b01010011: data1 <= -12'h117;
               8'b01010100: data1 <=  12'h0a3;
               8'b01010101: data1 <=  12'h302;
               8'b01010110: data1 <=  12'h13f;
               8'b01010111: data1 <=  12'h000;
               8'b01011000: data1 <=  12'h15c;
               8'b01011001: data1 <=  12'h024;
               8'b01011010: data1 <=  12'h024;
               8'b01011011: data1 <= -12'h060;
               8'b01011100: data1 <=  12'h01c;
               8'b01011101: data1 <=  12'h08a;
               8'b01011110: data1 <= -12'h00d;
               8'b01011111: data1 <=  12'h077;
               8'b01100000: data1 <= -12'h022;
               8'b01100001: data1 <= -12'h02c;
               8'b01100010: data1 <= -12'h064;
               8'b01100011: data1 <=  12'h00f;
               8'b01100100: data1 <= -12'h032;
               8'b01100101: data1 <= -12'h013;
               8'b01100110: data1 <=  12'h13a;
               8'b01100111: data1 <=  12'h075;
               8'b01101000: data1 <=  12'h050;
               8'b01101001: data1 <= -12'h077;
               8'b01101010: data1 <= -12'h077;
               8'b01101011: data1 <=  12'h050;
               8'b01101100: data1 <=  12'h011;
               8'b01101101: data1 <= -12'h091;
               8'b01101110: data1 <= -12'h042;
               8'b01101111: data1 <= -12'h05a;
               8'b01110000: data1 <= -12'h05d;
               8'b01110001: data1 <=  12'h044;
               8'b01110010: data1 <= -12'h036;
               8'b01110011: data1 <= -12'h08a;
               8'b01110100: data1 <=  12'h045;
               8'b01110101: data1 <=  12'h00d;
               8'b01110110: data1 <=  12'h156;
               8'b01110111: data1 <=  12'h420;
               8'b01111000: data1 <= -12'h095;
               8'b01111001: data1 <= -12'h043;
               8'b01111010: data1 <= -12'h00f;
               8'b01111011: data1 <= -12'h01a;
               8'b01111100: data1 <= -12'h00f;
               8'b01111101: data1 <= -12'h0ba;
               8'b01111110: data1 <= -12'h062;
               8'b01111111: data1 <= -12'h13d;
               8'b10000000: data1 <=  12'h060;
               8'b10000001: data1 <= -12'h00a;
               8'b10000010: data1 <=  12'h1eb;
               8'b10000011: data1 <=  12'h009;
               8'b10000100: data1 <=  12'h11d;
               8'b10000101: data1 <= -12'h0bf;
               8'b10000110: data1 <= -12'h0cd;
               8'b10000111: data1 <=  12'h07b;
               default: data1 <= 0;
           endcase
        end

endmodule: featureThreshold_rom
