module failVal_rom
  #(
     parameter W_DATA = 13,
     parameter W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1

     );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               12'b000000000000: data1 <= 13'h0216;
               12'b000000000001: data1 <= -13'h01dd;
               12'b000000000010: data1 <= -13'h0182;
               12'b000000000011: data1 <= -13'h00df;
               12'b000000000100: data1 <= -13'h00c7;
               12'b000000000101: data1 <= 13'h008e;
               12'b000000000110: data1 <= -13'h01b0;
               12'b000000000111: data1 <= -13'h017a;
               12'b000000001000: data1 <= -13'h00db;
               12'b000000001001: data1 <= 13'h013e;
               12'b000000001010: data1 <= -13'h019e;
               12'b000000001011: data1 <= -13'h01f1;
               12'b000000001100: data1 <= -13'h008e;
               12'b000000001101: data1 <= 13'h0044;
               12'b000000001110: data1 <= -13'h02ac;
               12'b000000001111: data1 <= -13'h0115;
               12'b000000010000: data1 <= -13'h005a;
               12'b000000010001: data1 <= 13'h00ed;
               12'b000000010010: data1 <= 13'h0128;
               12'b000000010011: data1 <= -13'h006b;
               12'b000000010100: data1 <= 13'h0175;
               12'b000000010101: data1 <= 13'h011e;
               12'b000000010110: data1 <= -13'h0059;
               12'b000000010111: data1 <= -13'h009b;
               12'b000000011000: data1 <= 13'h0063;
               12'b000000011001: data1 <= -13'h0103;
               12'b000000011010: data1 <= -13'h01a5;
               12'b000000011011: data1 <= 13'h0076;
               12'b000000011100: data1 <= -13'h00a7;
               12'b000000011101: data1 <= -13'h0165;
               12'b000000011110: data1 <= -13'h0081;
               12'b000000011111: data1 <= 13'h005d;
               12'b000000100000: data1 <= -13'h004d;
               12'b000000100001: data1 <= -13'h0067;
               12'b000000100010: data1 <= 13'h010d;
               12'b000000100011: data1 <= -13'h01a0;
               12'b000000100100: data1 <= 13'h0048;
               12'b000000100101: data1 <= -13'h0103;
               12'b000000100110: data1 <= -13'h002a;
               12'b000000100111: data1 <= 13'h0184;
               12'b000000101000: data1 <= 13'h01c3;
               12'b000000101001: data1 <= -13'h0050;
               12'b000000101010: data1 <= -13'h0019;
               12'b000000101011: data1 <= -13'h0067;
               12'b000000101100: data1 <= 13'h002b;
               12'b000000101101: data1 <= 13'h00e3;
               12'b000000101110: data1 <= -13'h005f;
               12'b000000101111: data1 <= 13'h0010;
               12'b000000110000: data1 <= -13'h01bf;
               12'b000000110001: data1 <= -13'h00f0;
               12'b000000110010: data1 <= -13'h000d;
               12'b000000110011: data1 <= -13'h01d4;

endmodule: failVal_rom
