module rect2_rom
  #(
     parameter W_DATA = 20,
     parameter W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );
     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               8'b00000000: data1 <=  20'h00000;
               8'b00000001: data1 <=  20'h00000;
               8'b00000010: data1 <=  20'h00000;
               8'b00000011: data1 <=  20'h00000;
               8'b00000100: data1 <=  20'h00000;
               8'b00000101: data1 <=  20'h00000;
               8'b00000110: data1 <=  20'h00000;
               8'b00000111: data1 <=  20'h00000;
               8'b00001000: data1 <=  20'h00000;
               8'b00001001: data1 <=  20'h00000;
               8'b00001010: data1 <=  20'h00000;
               8'b00001011: data1 <=  20'h00000;
               8'b00001100: data1 <=  20'h00000;
               8'b00001101: data1 <=  20'h00000;
               8'b00001110: data1 <=  20'h00000;
               8'b00001111: data1 <=  20'h00000;
               8'b00010000: data1 <=  20'h00000;
               8'b00010001: data1 <=  20'h00000;
               8'b00010010: data1 <=  20'h00000;
               8'b00010011: data1 <=  20'h00000;
               8'b00010100: data1 <=  20'h00000;
               8'b00010101: data1 <=  20'h00000;
               8'b00010110: data1 <=  20'h00000;
               8'b00010111: data1 <=  20'h00000;
               8'b00011000: data1 <=  20'h00000;
               8'b00011001: data1 <=  20'h00000;
               8'b00011010: data1 <=  20'h00000;
               8'b00011011: data1 <=  20'h00000;
               8'b00011100: data1 <=  20'h00000;
               8'b00011101: data1 <=  20'h00000;
               8'b00011110: data1 <=  20'h00000;
               8'b00011111: data1 <=  20'h00000;
               8'b00100000: data1 <=  20'h00000;
               8'b00100001: data1 <=  20'h00000;
               8'b00100010: data1 <=  20'h00000;
               8'b00100011: data1 <=  20'h4e0e6;
               8'b00100100: data1 <=  20'h00000;
               8'b00100101: data1 <=  20'h00000;
               8'b00100110: data1 <=  20'h00000;
               8'b00100111: data1 <=  20'h00000;
               8'b00101000: data1 <=  20'h00000;
               8'b00101001: data1 <=  20'h00000;
               8'b00101010: data1 <=  20'h00000;
               8'b00101011: data1 <=  20'h00000;
               8'b00101100: data1 <=  20'h00000;
               8'b00101101: data1 <=  20'h00000;
               8'b00101110: data1 <=  20'h00000;
               8'b00101111: data1 <=  20'h00000;
               8'b00110000: data1 <=  20'h4c4e7;
               8'b00110001: data1 <=  20'h00000;
               8'b00110010: data1 <=  20'h00000;
               8'b00110011: data1 <=  20'h00000;
               8'b00110100: data1 <=  20'h00000;
               8'b00110101: data1 <=  20'h00000;
               8'b00110110: data1 <=  20'h00000;
               8'b00110111: data1 <=  20'h00000;
               8'b00111000: data1 <=  20'h7f0c3;
               8'b00111001: data1 <=  20'h00000;
               8'b00111010: data1 <=  20'h00000;
               8'b00111011: data1 <=  20'h00000;
               8'b00111100: data1 <=  20'h00000;
               8'b00111101: data1 <=  20'h00000;
               8'b00111110: data1 <=  20'h60903;
               8'b00111111: data1 <=  20'h00000;
               8'b01000000: data1 <=  20'h00000;
               8'b01000001: data1 <=  20'h00000;
               8'b01000010: data1 <=  20'h00000;
               8'b01000011: data1 <=  20'h00000;
               8'b01000100: data1 <=  20'h00000;
               8'b01000101: data1 <=  20'h00000;
               8'b01000110: data1 <=  20'h4dd47;
               8'b01000111: data1 <=  20'h00000;
               8'b01001000: data1 <=  20'h00000;
               8'b01001001: data1 <=  20'h00000;
               8'b01001010: data1 <=  20'h00000;
               8'b01001011: data1 <=  20'h47885;
               8'b01001100: data1 <=  20'h4e0e7;
               8'b01001101: data1 <=  20'h00000;
               8'b01001110: data1 <=  20'h00000;
               8'b01001111: data1 <=  20'h00000;
               8'b01010000: data1 <=  20'h00000;
               8'b01010001: data1 <=  20'h00000;
               8'b01010010: data1 <=  20'h00000;
               8'b01010011: data1 <=  20'h00000;
               8'b01010100: data1 <=  20'h00000;
               8'b01010101: data1 <=  20'h00000;
               8'b01010110: data1 <=  20'h00000;
               8'b01010111: data1 <=  20'h00000;
               8'b01011000: data1 <=  20'h00000;
               8'b01011001: data1 <=  20'h00000;
               8'b01011010: data1 <=  20'h00000;
               8'b01011011: data1 <=  20'h00000;
               8'b01011100: data1 <=  20'h00000;
               8'b01011101: data1 <=  20'h00000;
               8'b01011110: data1 <=  20'h00000;
               8'b01011111: data1 <=  20'h00000;
               8'b01100000: data1 <=  20'h00000;
               8'b01100001: data1 <=  20'h00000;
               8'b01100010: data1 <=  20'h00000;
               8'b01100011: data1 <=  20'h00000;
               8'b01100100: data1 <=  20'h00000;
               8'b01100101: data1 <=  20'h00000;
               8'b01100110: data1 <=  20'h00000;
               8'b01100111: data1 <=  20'h00000;
               8'b01101000: data1 <=  20'h00000;
               8'b01101001: data1 <=  20'h77543;
               8'b01101010: data1 <=  20'h00000;
               8'b01101011: data1 <=  20'h00000;
               8'b01101100: data1 <=  20'h00000;
               8'b01101101: data1 <=  20'h478c3;
               8'b01101110: data1 <=  20'h464c3;
               8'b01101111: data1 <=  20'h00000;
               8'b01110000: data1 <=  20'h00000;
               8'b01110001: data1 <=  20'h00000;
               8'b01110010: data1 <=  20'h00000;
               8'b01110011: data1 <=  20'h00000;
               8'b01110100: data1 <=  20'h00000;
               8'b01110101: data1 <=  20'h00000;
               8'b01110110: data1 <=  20'h60926;
               8'b01110111: data1 <=  20'h00000;
               8'b01111000: data1 <=  20'h47ce5;
               8'b01111001: data1 <=  20'h470a6;
               8'b01111010: data1 <=  20'h474c6;
               8'b01111011: data1 <=  20'h00000;
               8'b01111100: data1 <=  20'h00000;
               8'b01111101: data1 <=  20'h00000;
               8'b01111110: data1 <=  20'h00000;
               8'b01111111: data1 <=  20'h00000;
               8'b10000000: data1 <=  20'h00000;
               8'b10000001: data1 <=  20'h00000;
               8'b10000010: data1 <=  20'h00000;
               8'b10000011: data1 <=  20'h00000;
               8'b10000100: data1 <=  20'h00000;
               8'b10000101: data1 <=  20'h00000;
               8'b10000110: data1 <=  20'h00000;
               8'b10000111: data1 <=  20'h00000;
               default: data1 <= 0;
           endcase
        end

endmodule: rect2_rom
