module weights1_rom
  #(
     parameter W_DATA = 3,
     parameter W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1

     );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               12'b000000000000: data1 <= 3'h3;
               12'b000000000001: data1 <= 3'h3;
               12'b000000000010: data1 <= 3'h3;
               12'b000000000011: data1 <= 3'h3;
               12'b000000000100: data1 <= 3'h2;
               12'b000000000101: data1 <= 3'h2;
               12'b000000000110: data1 <= 3'h2;
               12'b000000000111: data1 <= 3'h2;
               12'b000000001000: data1 <= 3'h2;
               12'b000000001001: data1 <= 3'h3;
               12'b000000001010: data1 <= 3'h3;
               12'b000000001011: data1 <= 3'h3;
               12'b000000001100: data1 <= 3'h3;
               12'b000000001101: data1 <= 3'h3;
               12'b000000001110: data1 <= 3'h2;
               12'b000000001111: data1 <= 3'h3;
               12'b000000010000: data1 <= 3'h3;
               12'b000000010001: data1 <= 3'h3;
               12'b000000010010: data1 <= 3'h3;
               12'b000000010011: data1 <= 3'h2;
               12'b000000010100: data1 <= 3'h3;
               12'b000000010101: data1 <= 3'h3;
               12'b000000010110: data1 <= 3'h3;
               12'b000000010111: data1 <= 3'h3;
               12'b000000011000: data1 <= 3'h2;
               12'b000000011001: data1 <= 3'h3;
               12'b000000011010: data1 <= 3'h2;
               12'b000000011011: data1 <= 3'h2;
               12'b000000011100: data1 <= 3'h3;
               12'b000000011101: data1 <= 3'h2;
               12'b000000011110: data1 <= 3'h3;
               12'b000000011111: data1 <= 3'h3;
               12'b000000100000: data1 <= 3'h2;
               12'b000000100001: data1 <= 3'h2;
               12'b000000100010: data1 <= 3'h3;
               12'b000000100011: data1 <= 3'h2;
               12'b000000100100: data1 <= 3'h3;
               12'b000000100101: data1 <= 3'h2;
               12'b000000100110: data1 <= 3'h2;
               12'b000000100111: data1 <= 3'h3;
               12'b000000101000: data1 <= 3'h2;
               12'b000000101001: data1 <= 3'h2;
               12'b000000101010: data1 <= 3'h3;
               12'b000000101011: data1 <= 3'h3;
               12'b000000101100: data1 <= 3'h2;
               12'b000000101101: data1 <= 3'h3;
               12'b000000101110: data1 <= 3'h2;
               12'b000000101111: data1 <= 3'h2;
               12'b000000110000: data1 <= 3'h2;
               12'b000000110001: data1 <= 3'h2;
               12'b000000110010: data1 <= 3'h2;
               12'b000000110011: data1 <= 3'h3;
               default: data1 <= 0;
           endcase
        end

endmodule: weights1_rom
