module rect1_rom
  #(
     parameter W_DATA = 20,
     parameter W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );
     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               8'b00000000: data1 <=  20'h2d583;
               8'b00000001: data1 <=  20'h1b887;
               8'b00000010: data1 <=  20'h4be43;
               8'b00000011: data1 <=  20'h7f122;
               8'b00000100: data1 <=  20'h20853;
               8'b00000101: data1 <=  20'h52d88;
               8'b00000110: data1 <=  20'h46183;
               8'b00000111: data1 <=  20'h79885;
               8'b00001000: data1 <=  20'h13ce3;
               8'b00001001: data1 <=  20'h33982;
               8'b00001010: data1 <=  20'h1b887;
               8'b00001011: data1 <=  20'h4b664;
               8'b00001100: data1 <=  20'h0e903;
               8'b00001101: data1 <=  20'h59cc5;
               8'b00001110: data1 <=  20'h461c5;
               8'b00001111: data1 <=  20'h141c3;
               8'b00010000: data1 <=  20'h48c66;
               8'b00010001: data1 <=  20'h2184a;
               8'b00010010: data1 <=  20'h3504a;
               8'b00010011: data1 <=  20'h20449;
               8'b00010100: data1 <=  20'h0504b;
               8'b00010101: data1 <=  20'h2790d;
               8'b00010110: data1 <=  20'h28449;
               8'b00010111: data1 <=  20'h7ed42;
               8'b00011000: data1 <=  20'h529c6;
               8'b00011001: data1 <=  20'h14d03;
               8'b00011010: data1 <=  20'h461e3;
               8'b00011011: data1 <=  20'h538a7;
               8'b00011100: data1 <=  20'h2204a;
               8'b00011101: data1 <=  20'h4c866;
               8'b00011110: data1 <=  20'h858c3;
               8'b00011111: data1 <=  20'h335a2;
               8'b00100000: data1 <=  20'h0ac6f;
               8'b00100001: data1 <=  20'h0746f;
               8'b00100010: data1 <=  20'h3410f;
               8'b00100011: data1 <=  20'h26ce6;
               8'b00100100: data1 <=  20'h64aa4;
               8'b00100101: data1 <=  20'h08c4a;
               8'b00100110: data1 <=  20'h51d4a;
               8'b00100111: data1 <=  20'h06c4d;
               8'b00101000: data1 <=  20'h1184d;
               8'b00101001: data1 <=  20'h22173;
               8'b00101010: data1 <=  20'h1e049;
               8'b00101011: data1 <=  20'h1344b;
               8'b00101100: data1 <=  20'h09449;
               8'b00101101: data1 <=  20'h2be61;
               8'b00101110: data1 <=  20'h09449;
               8'b00101111: data1 <=  20'h08c49;
               8'b00110000: data1 <=  20'h224e7;
               8'b00110001: data1 <=  20'h45241;
               8'b00110010: data1 <=  20'h5584b;
               8'b00110011: data1 <=  20'h2bcc3;
               8'b00110100: data1 <=  20'h2d583;
               8'b00110101: data1 <=  20'h21c86;
               8'b00110110: data1 <=  20'h08505;
               8'b00110111: data1 <=  20'h4c242;
               8'b00111000: data1 <=  20'h6acc3;
               8'b00111001: data1 <=  20'h1784d;
               8'b00111010: data1 <=  20'h1384d;
               8'b00111011: data1 <=  20'h08517;
               8'b00111100: data1 <=  20'h45104;
               8'b00111101: data1 <=  20'h5b067;
               8'b00111110: data1 <=  20'h4bd03;
               8'b00111111: data1 <=  20'h33982;
               8'b01000000: data1 <=  20'h534c6;
               8'b01000001: data1 <=  20'h6e122;
               8'b01000010: data1 <=  20'h70e41;
               8'b01000011: data1 <=  20'h3fa06;
               8'b01000100: data1 <=  20'h06c54;
               8'b01000101: data1 <=  20'h07241;
               8'b01000110: data1 <=  20'h1f947;
               8'b01000111: data1 <=  20'h4c5c4;
               8'b01001000: data1 <=  20'h6b0e3;
               8'b01001001: data1 <=  20'h6dd22;
               8'b01001010: data1 <=  20'h6a922;
               8'b01001011: data1 <=  20'h29485;
               8'b01001100: data1 <=  20'h208e7;
               8'b01001101: data1 <=  20'h02885;
               8'b01001110: data1 <=  20'h150c3;
               8'b01001111: data1 <=  20'h28449;
               8'b01010000: data1 <=  20'h02449;
               8'b01010001: data1 <=  20'h28849;
               8'b01010010: data1 <=  20'h28049;
               8'b01010011: data1 <=  20'h344c4;
               8'b01010100: data1 <=  20'h14583;
               8'b01010101: data1 <=  20'h02106;
               8'b01010110: data1 <=  20'h45e04;
               8'b01010111: data1 <=  20'h28466;
               8'b01011000: data1 <=  20'h7f103;
               8'b01011001: data1 <=  20'h28449;
               8'b01011010: data1 <=  20'h538a4;
               8'b01011011: data1 <=  20'h28449;
               8'b01011100: data1 <=  20'h28449;
               8'b01011101: data1 <=  20'h72cc6;
               8'b01011110: data1 <=  20'h90241;
               8'b01011111: data1 <=  20'h4d885;
               8'b01100000: data1 <=  20'h4c905;
               8'b01100001: data1 <=  20'h33d42;
               8'b01100010: data1 <=  20'h64142;
               8'b01100011: data1 <=  20'h78641;
               8'b01100100: data1 <=  20'h0cec1;
               8'b01100101: data1 <=  20'h6be41;
               8'b01100110: data1 <=  20'h1a46f;
               8'b01100111: data1 <=  20'h1e04a;
               8'b01101000: data1 <=  20'h1984a;
               8'b01101001: data1 <=  20'h67143;
               8'b01101010: data1 <=  20'h4c089;
               8'b01101011: data1 <=  20'h03849;
               8'b01101100: data1 <=  20'h40866;
               8'b01101101: data1 <=  20'h364c3;
               8'b01101110: data1 <=  20'h320c3;
               8'b01101111: data1 <=  20'h03849;
               8'b01110000: data1 <=  20'h02049;
               8'b01110001: data1 <=  20'h66122;
               8'b01110010: data1 <=  20'h70922;
               8'b01110011: data1 <=  20'h3504a;
               8'b01110100: data1 <=  20'h790c3;
               8'b01110101: data1 <=  20'h45681;
               8'b01110110: data1 <=  20'h38d26;
               8'b01110111: data1 <=  20'h00d38;
               8'b01111000: data1 <=  20'h26ce5;
               8'b01111001: data1 <=  20'h22ca6;
               8'b01111010: data1 <=  20'h204c6;
               8'b01111011: data1 <=  20'h5ee41;
               8'b01111100: data1 <=  20'h6bd04;
               8'b01111101: data1 <=  20'h77a43;
               8'b01111110: data1 <=  20'h00c66;
               8'b01111111: data1 <=  20'h28092;
               8'b10000000: data1 <=  20'h0844e;
               8'b10000001: data1 <=  20'h13a61;
               8'b10000010: data1 <=  20'h3516d;
               8'b10000011: data1 <=  20'h46d62;
               8'b10000100: data1 <=  20'h4c4aa;
               8'b10000101: data1 <=  20'h68086;
               8'b10000110: data1 <=  20'h65086;
               8'b10000111: data1 <=  20'h240a4;
               default: data1 <= 0;
           endcase
        end

endmodule: rect1_rom
