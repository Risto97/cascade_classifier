module rect0_rom
  #(
     parameter W_DATA = 20,
     parameter W_ADDR = 8
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1
    );
     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               8'b00000000: data1 <=  20'h1a989;
               8'b00000001: data1 <=  20'h1a987;
               8'b00000010: data1 <=  20'h39249;
               8'b00000011: data1 <=  20'h72926;
               8'b00000100: data1 <=  20'h20093;
               8'b00000101: data1 <=  20'h20d90;
               8'b00000110: data1 <=  20'h33586;
               8'b00000111: data1 <=  20'h5a48a;
               8'b00001000: data1 <=  20'h010e6;
               8'b00001001: data1 <=  20'h27186;
               8'b00001010: data1 <=  20'h1a987;
               8'b00001011: data1 <=  20'h3266c;
               8'b00001100: data1 <=  20'h0cb03;
               8'b00001101: data1 <=  20'h3a8cf;
               8'b00001110: data1 <=  20'h26dca;
               8'b00001111: data1 <=  20'h015c9;
               8'b00010000: data1 <=  20'h48126;
               8'b00010001: data1 <=  20'h210ca;
               8'b00010010: data1 <=  20'h348ca;
               8'b00010011: data1 <=  20'h1fc89;
               8'b00010100: data1 <=  20'h048cb;
               8'b00010101: data1 <=  20'h25b0d;
               8'b00010110: data1 <=  20'h27cc9;
               8'b00010111: data1 <=  20'h72546;
               8'b00011000: data1 <=  20'h2d1cc;
               8'b00011001: data1 <=  20'h12f03;
               8'b00011010: data1 <=  20'h335e6;
               8'b00011011: data1 <=  20'h27cae;
               8'b00011100: data1 <=  20'h218ca;
               8'b00011101: data1 <=  20'h2706c;
               8'b00011110: data1 <=  20'h84243;
               8'b00011111: data1 <=  20'h26da6;
               8'b00100000: data1 <=  20'h0accf;
               8'b00100001: data1 <=  20'h068cf;
               8'b00100010: data1 <=  20'h3230f;
               8'b00100011: data1 <=  20'h26dcc;
               8'b00100100: data1 <=  20'h4baac;
               8'b00100101: data1 <=  20'h0848a;
               8'b00100110: data1 <=  20'h51e8a;
               8'b00100111: data1 <=  20'h064cd;
               8'b00101000: data1 <=  20'h1188d;
               8'b00101001: data1 <=  20'h1f6d3;
               8'b00101010: data1 <=  20'h1d8c9;
               8'b00101011: data1 <=  20'h12ccb;
               8'b00101100: data1 <=  20'h09489;
               8'b00101101: data1 <=  20'h25a63;
               8'b00101110: data1 <=  20'h09489;
               8'b00101111: data1 <=  20'h08489;
               8'b00110000: data1 <=  20'h209ce;
               8'b00110001: data1 <=  20'h3ee42;
               8'b00110010: data1 <=  20'h5588b;
               8'b00110011: data1 <=  20'h190c9;
               8'b00110100: data1 <=  20'h1a989;
               8'b00110101: data1 <=  20'h20d86;
               8'b00110110: data1 <=  20'h06705;
               8'b00110111: data1 <=  20'h3fa46;
               8'b00111000: data1 <=  20'h6ad86;
               8'b00111001: data1 <=  20'h1788d;
               8'b00111010: data1 <=  20'h1308d;
               8'b00111011: data1 <=  20'h06717;
               8'b00111100: data1 <=  20'h2c10c;
               8'b00111101: data1 <=  20'h2f46e;
               8'b00111110: data1 <=  20'h4be06;
               8'b00111111: data1 <=  20'h27186;
               8'b01000000: data1 <=  20'h2dccc;
               8'b01000001: data1 <=  20'h61926;
               8'b01000010: data1 <=  20'h6aa43;
               8'b01000011: data1 <=  20'h1a20c;
               8'b01000100: data1 <=  20'h06494;
               8'b01000101: data1 <=  20'h00e42;
               8'b01000110: data1 <=  20'h1fa8e;
               8'b01000111: data1 <=  20'h335cc;
               8'b01001000: data1 <=  20'h584e9;
               8'b01001001: data1 <=  20'h61526;
               8'b01001010: data1 <=  20'h5e126;
               8'b01001011: data1 <=  20'h2850a;
               8'b01001100: data1 <=  20'h209ce;
               8'b01001101: data1 <=  20'h01985;
               8'b01001110: data1 <=  20'h024c9;
               8'b01001111: data1 <=  20'h27cc9;
               8'b01010000: data1 <=  20'h01cc9;
               8'b01010001: data1 <=  20'h280c9;
               8'b01010010: data1 <=  20'h278c9;
               8'b01010011: data1 <=  20'h32e44;
               8'b01010100: data1 <=  20'h01989;
               8'b01010101: data1 <=  20'h00306;
               8'b01010110: data1 <=  20'h2ce0c;
               8'b01010111: data1 <=  20'h284c6;
               8'b01011000: data1 <=  20'h7d303;
               8'b01011001: data1 <=  20'h28489;
               8'b01011010: data1 <=  20'h525e4;
               8'b01011011: data1 <=  20'h28489;
               8'b01011100: data1 <=  20'h27c89;
               8'b01011101: data1 <=  20'h4d4cc;
               8'b01011110: data1 <=  20'h89e42;
               8'b01011111: data1 <=  20'h2e48a;
               8'b01100000: data1 <=  20'h2d50a;
               8'b01100001: data1 <=  20'h27546;
               8'b01100010: data1 <=  20'h57944;
               8'b01100011: data1 <=  20'h72242;
               8'b01100100: data1 <=  20'h06ac3;
               8'b01100101: data1 <=  20'h65a43;
               8'b01100110: data1 <=  20'h198cf;
               8'b01100111: data1 <=  20'h1e08a;
               8'b01101000: data1 <=  20'h1908a;
               8'b01101001: data1 <=  20'h64a86;
               8'b01101010: data1 <=  20'h4b109;
               8'b01101011: data1 <=  20'h030c9;
               8'b01101100: data1 <=  20'h3fcc6;
               8'b01101101: data1 <=  20'h34d86;
               8'b01101110: data1 <=  20'h32186;
               8'b01101111: data1 <=  20'h030c9;
               8'b01110000: data1 <=  20'h018c9;
               8'b01110001: data1 <=  20'h59926;
               8'b01110010: data1 <=  20'h64126;
               8'b01110011: data1 <=  20'h348ca;
               8'b01110100: data1 <=  20'h77983;
               8'b01110101: data1 <=  20'h3f282;
               8'b01110110: data1 <=  20'h38e4c;
               8'b01110111: data1 <=  20'h00e58;
               8'b01111000: data1 <=  20'h26dca;
               8'b01111001: data1 <=  20'h2194c;
               8'b01111010: data1 <=  20'h2058c;
               8'b01111011: data1 <=  20'h58a43;
               8'b01111100: data1 <=  20'h52d08;
               8'b01111101: data1 <=  20'h64e46;
               8'b01111110: data1 <=  20'h000c6;
               8'b01111111: data1 <=  20'h27192;
               8'b10000000: data1 <=  20'h07c8e;
               8'b10000001: data1 <=  20'h0d662;
               8'b10000010: data1 <=  20'h326cd;
               8'b10000011: data1 <=  20'h3a564;
               8'b10000100: data1 <=  20'h4b1ea;
               8'b10000101: data1 <=  20'h67186;
               8'b10000110: data1 <=  20'h64186;
               8'b10000111: data1 <=  20'h0b0ac;
               default: data1 <= 0;
           endcase
        end

endmodule: rect0_rom
