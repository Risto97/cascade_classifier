module weights0_rom
  #(
     W_DATA = 3,
     DEPTH = 2913,
     W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input ena,
     input [W_ADDR-1:0] addra,
     output [W_DATA-1:0] doa
    );

     logic [W_DATA-1:0] mem [DEPTH-1:0];

     always_ff @(posedge clk)
        begin
           if(ena)
              doa = mem[addra];
        end

     initial begin
         mem[0] = -3'h1;
         mem[1] = -3'h1;
         mem[2] = -3'h1;
         mem[3] = -3'h1;
         mem[4] = -3'h1;
         mem[5] = -3'h1;
         mem[6] = -3'h1;
         mem[7] = -3'h1;
         mem[8] = -3'h1;
         mem[9] = -3'h1;
         mem[10] = -3'h1;
         mem[11] = -3'h1;
         mem[12] = -3'h1;
         mem[13] = -3'h1;
         mem[14] = -3'h1;
         mem[15] = -3'h1;
         mem[16] = -3'h1;
         mem[17] = -3'h1;
         mem[18] = -3'h1;
         mem[19] = -3'h1;
         mem[20] = -3'h1;
         mem[21] = -3'h1;
         mem[22] = -3'h1;
         mem[23] = -3'h1;
         mem[24] = -3'h1;
         mem[25] = -3'h1;
         mem[26] = -3'h1;
         mem[27] = -3'h1;
         mem[28] = -3'h1;
         mem[29] = -3'h1;
         mem[30] = -3'h1;
         mem[31] = -3'h1;
         mem[32] = -3'h1;
         mem[33] = -3'h1;
         mem[34] = -3'h1;
         mem[35] = -3'h1;
         mem[36] = -3'h1;
         mem[37] = -3'h1;
         mem[38] = -3'h1;
         mem[39] = -3'h1;
         mem[40] = -3'h1;
         mem[41] = -3'h1;
         mem[42] = -3'h1;
         mem[43] = -3'h1;
         mem[44] = -3'h1;
         mem[45] = -3'h1;
         mem[46] = -3'h1;
         mem[47] = -3'h1;
         mem[48] = -3'h1;
         mem[49] = -3'h1;
         mem[50] = -3'h1;
         mem[51] = -3'h1;
         mem[52] = -3'h1;
         mem[53] = -3'h1;
         mem[54] = -3'h1;
         mem[55] = -3'h1;
         mem[56] = -3'h1;
         mem[57] = -3'h1;
         mem[58] = -3'h1;
         mem[59] = -3'h1;
         mem[60] = -3'h1;
         mem[61] = -3'h1;
         mem[62] = -3'h1;
         mem[63] = -3'h1;
         mem[64] = -3'h1;
         mem[65] = -3'h1;
         mem[66] = -3'h1;
         mem[67] = -3'h1;
         mem[68] = -3'h1;
         mem[69] = -3'h1;
         mem[70] = -3'h1;
         mem[71] = -3'h1;
         mem[72] = -3'h1;
         mem[73] = -3'h1;
         mem[74] = -3'h1;
         mem[75] = -3'h1;
         mem[76] = -3'h1;
         mem[77] = -3'h1;
         mem[78] = -3'h1;
         mem[79] = -3'h1;
         mem[80] = -3'h1;
         mem[81] = -3'h1;
         mem[82] = -3'h1;
         mem[83] = -3'h1;
         mem[84] = -3'h1;
         mem[85] = -3'h1;
         mem[86] = -3'h1;
         mem[87] = -3'h1;
         mem[88] = -3'h1;
         mem[89] = -3'h1;
         mem[90] = -3'h1;
         mem[91] = -3'h1;
         mem[92] = -3'h1;
         mem[93] = -3'h1;
         mem[94] = -3'h1;
         mem[95] = -3'h1;
         mem[96] = -3'h1;
         mem[97] = -3'h1;
         mem[98] = -3'h1;
         mem[99] = -3'h1;
         mem[100] = -3'h1;
         mem[101] = -3'h1;
         mem[102] = -3'h1;
         mem[103] = -3'h1;
         mem[104] = -3'h1;
         mem[105] = -3'h1;
         mem[106] = -3'h1;
         mem[107] = -3'h1;
         mem[108] = -3'h1;
         mem[109] = -3'h1;
         mem[110] = -3'h1;
         mem[111] = -3'h1;
         mem[112] = -3'h1;
         mem[113] = -3'h1;
         mem[114] = -3'h1;
         mem[115] = -3'h1;
         mem[116] = -3'h1;
         mem[117] = -3'h1;
         mem[118] = -3'h1;
         mem[119] = -3'h1;
         mem[120] = -3'h1;
         mem[121] = -3'h1;
         mem[122] = -3'h1;
         mem[123] = -3'h1;
         mem[124] = -3'h1;
         mem[125] = -3'h1;
         mem[126] = -3'h1;
         mem[127] = -3'h1;
         mem[128] = -3'h1;
         mem[129] = -3'h1;
         mem[130] = -3'h1;
         mem[131] = -3'h1;
         mem[132] = -3'h1;
         mem[133] = -3'h1;
         mem[134] = -3'h1;
         mem[135] = -3'h1;
         mem[136] = -3'h1;
         mem[137] = -3'h1;
         mem[138] = -3'h1;
         mem[139] = -3'h1;
         mem[140] = -3'h1;
         mem[141] = -3'h1;
         mem[142] = -3'h1;
         mem[143] = -3'h1;
         mem[144] = -3'h1;
         mem[145] = -3'h1;
         mem[146] = -3'h1;
         mem[147] = -3'h1;
         mem[148] = -3'h1;
         mem[149] = -3'h1;
         mem[150] = -3'h1;
         mem[151] = -3'h1;
         mem[152] = -3'h1;
         mem[153] = -3'h1;
         mem[154] = -3'h1;
         mem[155] = -3'h1;
         mem[156] = -3'h1;
         mem[157] = -3'h1;
         mem[158] = -3'h1;
         mem[159] = -3'h1;
         mem[160] = -3'h1;
         mem[161] = -3'h1;
         mem[162] = -3'h1;
         mem[163] = -3'h1;
         mem[164] = -3'h1;
         mem[165] = -3'h1;
         mem[166] = -3'h1;
         mem[167] = -3'h1;
         mem[168] = -3'h1;
         mem[169] = -3'h1;
         mem[170] = -3'h1;
         mem[171] = -3'h1;
         mem[172] = -3'h1;
         mem[173] = -3'h1;
         mem[174] = -3'h1;
         mem[175] = -3'h1;
         mem[176] = -3'h1;
         mem[177] = -3'h1;
         mem[178] = -3'h1;
         mem[179] = -3'h1;
         mem[180] = -3'h1;
         mem[181] = -3'h1;
         mem[182] = -3'h1;
         mem[183] = -3'h1;
         mem[184] = -3'h1;
         mem[185] = -3'h1;
         mem[186] = -3'h1;
         mem[187] = -3'h1;
         mem[188] = -3'h1;
         mem[189] = -3'h1;
         mem[190] = -3'h1;
         mem[191] = -3'h1;
         mem[192] = -3'h1;
         mem[193] = -3'h1;
         mem[194] = -3'h1;
         mem[195] = -3'h1;
         mem[196] = -3'h1;
         mem[197] = -3'h1;
         mem[198] = -3'h1;
         mem[199] = -3'h1;
         mem[200] = -3'h1;
         mem[201] = -3'h1;
         mem[202] = -3'h1;
         mem[203] = -3'h1;
         mem[204] = -3'h1;
         mem[205] = -3'h1;
         mem[206] = -3'h1;
         mem[207] = -3'h1;
         mem[208] = -3'h1;
         mem[209] = -3'h1;
         mem[210] = -3'h1;
         mem[211] = -3'h1;
         mem[212] = -3'h1;
         mem[213] = -3'h1;
         mem[214] = -3'h1;
         mem[215] = -3'h1;
         mem[216] = -3'h1;
         mem[217] = -3'h1;
         mem[218] = -3'h1;
         mem[219] = -3'h1;
         mem[220] = -3'h1;
         mem[221] = -3'h1;
         mem[222] = -3'h1;
         mem[223] = -3'h1;
         mem[224] = -3'h1;
         mem[225] = -3'h1;
         mem[226] = -3'h1;
         mem[227] = -3'h1;
         mem[228] = -3'h1;
         mem[229] = -3'h1;
         mem[230] = -3'h1;
         mem[231] = -3'h1;
         mem[232] = -3'h1;
         mem[233] = -3'h1;
         mem[234] = -3'h1;
         mem[235] = -3'h1;
         mem[236] = -3'h1;
         mem[237] = -3'h1;
         mem[238] = -3'h1;
         mem[239] = -3'h1;
         mem[240] = -3'h1;
         mem[241] = -3'h1;
         mem[242] = -3'h1;
         mem[243] = -3'h1;
         mem[244] = -3'h1;
         mem[245] = -3'h1;
         mem[246] = -3'h1;
         mem[247] = -3'h1;
         mem[248] = -3'h1;
         mem[249] = -3'h1;
         mem[250] = -3'h1;
         mem[251] = -3'h1;
         mem[252] = -3'h1;
         mem[253] = -3'h1;
         mem[254] = -3'h1;
         mem[255] = -3'h1;
         mem[256] = -3'h1;
         mem[257] = -3'h1;
         mem[258] = -3'h1;
         mem[259] = -3'h1;
         mem[260] = -3'h1;
         mem[261] = -3'h1;
         mem[262] = -3'h1;
         mem[263] = -3'h1;
         mem[264] = -3'h1;
         mem[265] = -3'h1;
         mem[266] = -3'h1;
         mem[267] = -3'h1;
         mem[268] = -3'h1;
         mem[269] = -3'h1;
         mem[270] = -3'h1;
         mem[271] = -3'h1;
         mem[272] = -3'h1;
         mem[273] = -3'h1;
         mem[274] = -3'h1;
         mem[275] = -3'h1;
         mem[276] = -3'h1;
         mem[277] = -3'h1;
         mem[278] = -3'h1;
         mem[279] = -3'h1;
         mem[280] = -3'h1;
         mem[281] = -3'h1;
         mem[282] = -3'h1;
         mem[283] = -3'h1;
         mem[284] = -3'h1;
         mem[285] = -3'h1;
         mem[286] = -3'h1;
         mem[287] = -3'h1;
         mem[288] = -3'h1;
         mem[289] = -3'h1;
         mem[290] = -3'h1;
         mem[291] = -3'h1;
         mem[292] = -3'h1;
         mem[293] = -3'h1;
         mem[294] = -3'h1;
         mem[295] = -3'h1;
         mem[296] = -3'h1;
         mem[297] = -3'h1;
         mem[298] = -3'h1;
         mem[299] = -3'h1;
         mem[300] = -3'h1;
         mem[301] = -3'h1;
         mem[302] = -3'h1;
         mem[303] = -3'h1;
         mem[304] = -3'h1;
         mem[305] = -3'h1;
         mem[306] = -3'h1;
         mem[307] = -3'h1;
         mem[308] = -3'h1;
         mem[309] = -3'h1;
         mem[310] = -3'h1;
         mem[311] = -3'h1;
         mem[312] = -3'h1;
         mem[313] = -3'h1;
         mem[314] = -3'h1;
         mem[315] = -3'h1;
         mem[316] = -3'h1;
         mem[317] = -3'h1;
         mem[318] = -3'h1;
         mem[319] = -3'h1;
         mem[320] = -3'h1;
         mem[321] = -3'h1;
         mem[322] = -3'h1;
         mem[323] = -3'h1;
         mem[324] = -3'h1;
         mem[325] = -3'h1;
         mem[326] = -3'h1;
         mem[327] = -3'h1;
         mem[328] = -3'h1;
         mem[329] = -3'h1;
         mem[330] = -3'h1;
         mem[331] = -3'h1;
         mem[332] = -3'h1;
         mem[333] = -3'h1;
         mem[334] = -3'h1;
         mem[335] = -3'h1;
         mem[336] = -3'h1;
         mem[337] = -3'h1;
         mem[338] = -3'h1;
         mem[339] = -3'h1;
         mem[340] = -3'h1;
         mem[341] = -3'h1;
         mem[342] = -3'h1;
         mem[343] = -3'h1;
         mem[344] = -3'h1;
         mem[345] = -3'h1;
         mem[346] = -3'h1;
         mem[347] = -3'h1;
         mem[348] = -3'h1;
         mem[349] = -3'h1;
         mem[350] = -3'h1;
         mem[351] = -3'h1;
         mem[352] = -3'h1;
         mem[353] = -3'h1;
         mem[354] = -3'h1;
         mem[355] = -3'h1;
         mem[356] = -3'h1;
         mem[357] = -3'h1;
         mem[358] = -3'h1;
         mem[359] = -3'h1;
         mem[360] = -3'h1;
         mem[361] = -3'h1;
         mem[362] = -3'h1;
         mem[363] = -3'h1;
         mem[364] = -3'h1;
         mem[365] = -3'h1;
         mem[366] = -3'h1;
         mem[367] = -3'h1;
         mem[368] = -3'h1;
         mem[369] = -3'h1;
         mem[370] = -3'h1;
         mem[371] = -3'h1;
         mem[372] = -3'h1;
         mem[373] = -3'h1;
         mem[374] = -3'h1;
         mem[375] = -3'h1;
         mem[376] = -3'h1;
         mem[377] = -3'h1;
         mem[378] = -3'h1;
         mem[379] = -3'h1;
         mem[380] = -3'h1;
         mem[381] = -3'h1;
         mem[382] = -3'h1;
         mem[383] = -3'h1;
         mem[384] = -3'h1;
         mem[385] = -3'h1;
         mem[386] = -3'h1;
         mem[387] = -3'h1;
         mem[388] = -3'h1;
         mem[389] = -3'h1;
         mem[390] = -3'h1;
         mem[391] = -3'h1;
         mem[392] = -3'h1;
         mem[393] = -3'h1;
         mem[394] = -3'h1;
         mem[395] = -3'h1;
         mem[396] = -3'h1;
         mem[397] = -3'h1;
         mem[398] = -3'h1;
         mem[399] = -3'h1;
         mem[400] = -3'h1;
         mem[401] = -3'h1;
         mem[402] = -3'h1;
         mem[403] = -3'h1;
         mem[404] = -3'h1;
         mem[405] = -3'h1;
         mem[406] = -3'h1;
         mem[407] = -3'h1;
         mem[408] = -3'h1;
         mem[409] = -3'h1;
         mem[410] = -3'h1;
         mem[411] = -3'h1;
         mem[412] = -3'h1;
         mem[413] = -3'h1;
         mem[414] = -3'h1;
         mem[415] = -3'h1;
         mem[416] = -3'h1;
         mem[417] = -3'h1;
         mem[418] = -3'h1;
         mem[419] = -3'h1;
         mem[420] = -3'h1;
         mem[421] = -3'h1;
         mem[422] = -3'h1;
         mem[423] = -3'h1;
         mem[424] = -3'h1;
         mem[425] = -3'h1;
         mem[426] = -3'h1;
         mem[427] = -3'h1;
         mem[428] = -3'h1;
         mem[429] = -3'h1;
         mem[430] = -3'h1;
         mem[431] = -3'h1;
         mem[432] = -3'h1;
         mem[433] = -3'h1;
         mem[434] = -3'h1;
         mem[435] = -3'h1;
         mem[436] = -3'h1;
         mem[437] = -3'h1;
         mem[438] = -3'h1;
         mem[439] = -3'h1;
         mem[440] = -3'h1;
         mem[441] = -3'h1;
         mem[442] = -3'h1;
         mem[443] = -3'h1;
         mem[444] = -3'h1;
         mem[445] = -3'h1;
         mem[446] = -3'h1;
         mem[447] = -3'h1;
         mem[448] = -3'h1;
         mem[449] = -3'h1;
         mem[450] = -3'h1;
         mem[451] = -3'h1;
         mem[452] = -3'h1;
         mem[453] = -3'h1;
         mem[454] = -3'h1;
         mem[455] = -3'h1;
         mem[456] = -3'h1;
         mem[457] = -3'h1;
         mem[458] = -3'h1;
         mem[459] = -3'h1;
         mem[460] = -3'h1;
         mem[461] = -3'h1;
         mem[462] = -3'h1;
         mem[463] = -3'h1;
         mem[464] = -3'h1;
         mem[465] = -3'h1;
         mem[466] = -3'h1;
         mem[467] = -3'h1;
         mem[468] = -3'h1;
         mem[469] = -3'h1;
         mem[470] = -3'h1;
         mem[471] = -3'h1;
         mem[472] = -3'h1;
         mem[473] = -3'h1;
         mem[474] = -3'h1;
         mem[475] = -3'h1;
         mem[476] = -3'h1;
         mem[477] = -3'h1;
         mem[478] = -3'h1;
         mem[479] = -3'h1;
         mem[480] = -3'h1;
         mem[481] = -3'h1;
         mem[482] = -3'h1;
         mem[483] = -3'h1;
         mem[484] = -3'h1;
         mem[485] = -3'h1;
         mem[486] = -3'h1;
         mem[487] = -3'h1;
         mem[488] = -3'h1;
         mem[489] = -3'h1;
         mem[490] = -3'h1;
         mem[491] = -3'h1;
         mem[492] = -3'h1;
         mem[493] = -3'h1;
         mem[494] = -3'h1;
         mem[495] = -3'h1;
         mem[496] = -3'h1;
         mem[497] = -3'h1;
         mem[498] = -3'h1;
         mem[499] = -3'h1;
         mem[500] = -3'h1;
         mem[501] = -3'h1;
         mem[502] = -3'h1;
         mem[503] = -3'h1;
         mem[504] = -3'h1;
         mem[505] = -3'h1;
         mem[506] = -3'h1;
         mem[507] = -3'h1;
         mem[508] = -3'h1;
         mem[509] = -3'h1;
         mem[510] = -3'h1;
         mem[511] = -3'h1;
         mem[512] = -3'h1;
         mem[513] = -3'h1;
         mem[514] = -3'h1;
         mem[515] = -3'h1;
         mem[516] = -3'h1;
         mem[517] = -3'h1;
         mem[518] = -3'h1;
         mem[519] = -3'h1;
         mem[520] = -3'h1;
         mem[521] = -3'h1;
         mem[522] = -3'h1;
         mem[523] = -3'h1;
         mem[524] = -3'h1;
         mem[525] = -3'h1;
         mem[526] = -3'h1;
         mem[527] = -3'h1;
         mem[528] = -3'h1;
         mem[529] = -3'h1;
         mem[530] = -3'h1;
         mem[531] = -3'h1;
         mem[532] = -3'h1;
         mem[533] = -3'h1;
         mem[534] = -3'h1;
         mem[535] = -3'h1;
         mem[536] = -3'h1;
         mem[537] = -3'h1;
         mem[538] = -3'h1;
         mem[539] = -3'h1;
         mem[540] = -3'h1;
         mem[541] = -3'h1;
         mem[542] = -3'h1;
         mem[543] = -3'h1;
         mem[544] = -3'h1;
         mem[545] = -3'h1;
         mem[546] = -3'h1;
         mem[547] = -3'h1;
         mem[548] = -3'h1;
         mem[549] = -3'h1;
         mem[550] = -3'h1;
         mem[551] = -3'h1;
         mem[552] = -3'h1;
         mem[553] = -3'h1;
         mem[554] = -3'h1;
         mem[555] = -3'h1;
         mem[556] = -3'h1;
         mem[557] = -3'h1;
         mem[558] = -3'h1;
         mem[559] = -3'h1;
         mem[560] = -3'h1;
         mem[561] = -3'h1;
         mem[562] = -3'h1;
         mem[563] = -3'h1;
         mem[564] = -3'h1;
         mem[565] = -3'h1;
         mem[566] = -3'h1;
         mem[567] = -3'h1;
         mem[568] = -3'h1;
         mem[569] = -3'h1;
         mem[570] = -3'h1;
         mem[571] = -3'h1;
         mem[572] = -3'h1;
         mem[573] = -3'h1;
         mem[574] = -3'h1;
         mem[575] = -3'h1;
         mem[576] = -3'h1;
         mem[577] = -3'h1;
         mem[578] = -3'h1;
         mem[579] = -3'h1;
         mem[580] = -3'h1;
         mem[581] = -3'h1;
         mem[582] = -3'h1;
         mem[583] = -3'h1;
         mem[584] = -3'h1;
         mem[585] = -3'h1;
         mem[586] = -3'h1;
         mem[587] = -3'h1;
         mem[588] = -3'h1;
         mem[589] = -3'h1;
         mem[590] = -3'h1;
         mem[591] = -3'h1;
         mem[592] = -3'h1;
         mem[593] = -3'h1;
         mem[594] = -3'h1;
         mem[595] = -3'h1;
         mem[596] = -3'h1;
         mem[597] = -3'h1;
         mem[598] = -3'h1;
         mem[599] = -3'h1;
         mem[600] = -3'h1;
         mem[601] = -3'h1;
         mem[602] = -3'h1;
         mem[603] = -3'h1;
         mem[604] = -3'h1;
         mem[605] = -3'h1;
         mem[606] = -3'h1;
         mem[607] = -3'h1;
         mem[608] = -3'h1;
         mem[609] = -3'h1;
         mem[610] = -3'h1;
         mem[611] = -3'h1;
         mem[612] = -3'h1;
         mem[613] = -3'h1;
         mem[614] = -3'h1;
         mem[615] = -3'h1;
         mem[616] = -3'h1;
         mem[617] = -3'h1;
         mem[618] = -3'h1;
         mem[619] = -3'h1;
         mem[620] = -3'h1;
         mem[621] = -3'h1;
         mem[622] = -3'h1;
         mem[623] = -3'h1;
         mem[624] = -3'h1;
         mem[625] = -3'h1;
         mem[626] = -3'h1;
         mem[627] = -3'h1;
         mem[628] = -3'h1;
         mem[629] = -3'h1;
         mem[630] = -3'h1;
         mem[631] = -3'h1;
         mem[632] = -3'h1;
         mem[633] = -3'h1;
         mem[634] = -3'h1;
         mem[635] = -3'h1;
         mem[636] = -3'h1;
         mem[637] = -3'h1;
         mem[638] = -3'h1;
         mem[639] = -3'h1;
         mem[640] = -3'h1;
         mem[641] = -3'h1;
         mem[642] = -3'h1;
         mem[643] = -3'h1;
         mem[644] = -3'h1;
         mem[645] = -3'h1;
         mem[646] = -3'h1;
         mem[647] = -3'h1;
         mem[648] = -3'h1;
         mem[649] = -3'h1;
         mem[650] = -3'h1;
         mem[651] = -3'h1;
         mem[652] = -3'h1;
         mem[653] = -3'h1;
         mem[654] = -3'h1;
         mem[655] = -3'h1;
         mem[656] = -3'h1;
         mem[657] = -3'h1;
         mem[658] = -3'h1;
         mem[659] = -3'h1;
         mem[660] = -3'h1;
         mem[661] = -3'h1;
         mem[662] = -3'h1;
         mem[663] = -3'h1;
         mem[664] = -3'h1;
         mem[665] = -3'h1;
         mem[666] = -3'h1;
         mem[667] = -3'h1;
         mem[668] = -3'h1;
         mem[669] = -3'h1;
         mem[670] = -3'h1;
         mem[671] = -3'h1;
         mem[672] = -3'h1;
         mem[673] = -3'h1;
         mem[674] = -3'h1;
         mem[675] = -3'h1;
         mem[676] = -3'h1;
         mem[677] = -3'h1;
         mem[678] = -3'h1;
         mem[679] = -3'h1;
         mem[680] = -3'h1;
         mem[681] = -3'h1;
         mem[682] = -3'h1;
         mem[683] = -3'h1;
         mem[684] = -3'h1;
         mem[685] = -3'h1;
         mem[686] = -3'h1;
         mem[687] = -3'h1;
         mem[688] = -3'h1;
         mem[689] = -3'h1;
         mem[690] = -3'h1;
         mem[691] = -3'h1;
         mem[692] = -3'h1;
         mem[693] = -3'h1;
         mem[694] = -3'h1;
         mem[695] = -3'h1;
         mem[696] = -3'h1;
         mem[697] = -3'h1;
         mem[698] = -3'h1;
         mem[699] = -3'h1;
         mem[700] = -3'h1;
         mem[701] = -3'h1;
         mem[702] = -3'h1;
         mem[703] = -3'h1;
         mem[704] = -3'h1;
         mem[705] = -3'h1;
         mem[706] = -3'h1;
         mem[707] = -3'h1;
         mem[708] = -3'h1;
         mem[709] = -3'h1;
         mem[710] = -3'h1;
         mem[711] = -3'h1;
         mem[712] = -3'h1;
         mem[713] = -3'h1;
         mem[714] = -3'h1;
         mem[715] = -3'h1;
         mem[716] = -3'h1;
         mem[717] = -3'h1;
         mem[718] = -3'h1;
         mem[719] = -3'h1;
         mem[720] = -3'h1;
         mem[721] = -3'h1;
         mem[722] = -3'h1;
         mem[723] = -3'h1;
         mem[724] = -3'h1;
         mem[725] = -3'h1;
         mem[726] = -3'h1;
         mem[727] = -3'h1;
         mem[728] = -3'h1;
         mem[729] = -3'h1;
         mem[730] = -3'h1;
         mem[731] = -3'h1;
         mem[732] = -3'h1;
         mem[733] = -3'h1;
         mem[734] = -3'h1;
         mem[735] = -3'h1;
         mem[736] = -3'h1;
         mem[737] = -3'h1;
         mem[738] = -3'h1;
         mem[739] = -3'h1;
         mem[740] = -3'h1;
         mem[741] = -3'h1;
         mem[742] = -3'h1;
         mem[743] = -3'h1;
         mem[744] = -3'h1;
         mem[745] = -3'h1;
         mem[746] = -3'h1;
         mem[747] = -3'h1;
         mem[748] = -3'h1;
         mem[749] = -3'h1;
         mem[750] = -3'h1;
         mem[751] = -3'h1;
         mem[752] = -3'h1;
         mem[753] = -3'h1;
         mem[754] = -3'h1;
         mem[755] = -3'h1;
         mem[756] = -3'h1;
         mem[757] = -3'h1;
         mem[758] = -3'h1;
         mem[759] = -3'h1;
         mem[760] = -3'h1;
         mem[761] = -3'h1;
         mem[762] = -3'h1;
         mem[763] = -3'h1;
         mem[764] = -3'h1;
         mem[765] = -3'h1;
         mem[766] = -3'h1;
         mem[767] = -3'h1;
         mem[768] = -3'h1;
         mem[769] = -3'h1;
         mem[770] = -3'h1;
         mem[771] = -3'h1;
         mem[772] = -3'h1;
         mem[773] = -3'h1;
         mem[774] = -3'h1;
         mem[775] = -3'h1;
         mem[776] = -3'h1;
         mem[777] = -3'h1;
         mem[778] = -3'h1;
         mem[779] = -3'h1;
         mem[780] = -3'h1;
         mem[781] = -3'h1;
         mem[782] = -3'h1;
         mem[783] = -3'h1;
         mem[784] = -3'h1;
         mem[785] = -3'h1;
         mem[786] = -3'h1;
         mem[787] = -3'h1;
         mem[788] = -3'h1;
         mem[789] = -3'h1;
         mem[790] = -3'h1;
         mem[791] = -3'h1;
         mem[792] = -3'h1;
         mem[793] = -3'h1;
         mem[794] = -3'h1;
         mem[795] = -3'h1;
         mem[796] = -3'h1;
         mem[797] = -3'h1;
         mem[798] = -3'h1;
         mem[799] = -3'h1;
         mem[800] = -3'h1;
         mem[801] = -3'h1;
         mem[802] = -3'h1;
         mem[803] = -3'h1;
         mem[804] = -3'h1;
         mem[805] = -3'h1;
         mem[806] = -3'h1;
         mem[807] = -3'h1;
         mem[808] = -3'h1;
         mem[809] = -3'h1;
         mem[810] = -3'h1;
         mem[811] = -3'h1;
         mem[812] = -3'h1;
         mem[813] = -3'h1;
         mem[814] = -3'h1;
         mem[815] = -3'h1;
         mem[816] = -3'h1;
         mem[817] = -3'h1;
         mem[818] = -3'h1;
         mem[819] = -3'h1;
         mem[820] = -3'h1;
         mem[821] = -3'h1;
         mem[822] = -3'h1;
         mem[823] = -3'h1;
         mem[824] = -3'h1;
         mem[825] = -3'h1;
         mem[826] = -3'h1;
         mem[827] = -3'h1;
         mem[828] = -3'h1;
         mem[829] = -3'h1;
         mem[830] = -3'h1;
         mem[831] = -3'h1;
         mem[832] = -3'h1;
         mem[833] = -3'h1;
         mem[834] = -3'h1;
         mem[835] = -3'h1;
         mem[836] = -3'h1;
         mem[837] = -3'h1;
         mem[838] = -3'h1;
         mem[839] = -3'h1;
         mem[840] = -3'h1;
         mem[841] = -3'h1;
         mem[842] = -3'h1;
         mem[843] = -3'h1;
         mem[844] = -3'h1;
         mem[845] = -3'h1;
         mem[846] = -3'h1;
         mem[847] = -3'h1;
         mem[848] = -3'h1;
         mem[849] = -3'h1;
         mem[850] = -3'h1;
         mem[851] = -3'h1;
         mem[852] = -3'h1;
         mem[853] = -3'h1;
         mem[854] = -3'h1;
         mem[855] = -3'h1;
         mem[856] = -3'h1;
         mem[857] = -3'h1;
         mem[858] = -3'h1;
         mem[859] = -3'h1;
         mem[860] = -3'h1;
         mem[861] = -3'h1;
         mem[862] = -3'h1;
         mem[863] = -3'h1;
         mem[864] = -3'h1;
         mem[865] = -3'h1;
         mem[866] = -3'h1;
         mem[867] = -3'h1;
         mem[868] = -3'h1;
         mem[869] = -3'h1;
         mem[870] = -3'h1;
         mem[871] = -3'h1;
         mem[872] = -3'h1;
         mem[873] = -3'h1;
         mem[874] = -3'h1;
         mem[875] = -3'h1;
         mem[876] = -3'h1;
         mem[877] = -3'h1;
         mem[878] = -3'h1;
         mem[879] = -3'h1;
         mem[880] = -3'h1;
         mem[881] = -3'h1;
         mem[882] = -3'h1;
         mem[883] = -3'h1;
         mem[884] = -3'h1;
         mem[885] = -3'h1;
         mem[886] = -3'h1;
         mem[887] = -3'h1;
         mem[888] = -3'h1;
         mem[889] = -3'h1;
         mem[890] = -3'h1;
         mem[891] = -3'h1;
         mem[892] = -3'h1;
         mem[893] = -3'h1;
         mem[894] = -3'h1;
         mem[895] = -3'h1;
         mem[896] = -3'h1;
         mem[897] = -3'h1;
         mem[898] = -3'h1;
         mem[899] = -3'h1;
         mem[900] = -3'h1;
         mem[901] = -3'h1;
         mem[902] = -3'h1;
         mem[903] = -3'h1;
         mem[904] = -3'h1;
         mem[905] = -3'h1;
         mem[906] = -3'h1;
         mem[907] = -3'h1;
         mem[908] = -3'h1;
         mem[909] = -3'h1;
         mem[910] = -3'h1;
         mem[911] = -3'h1;
         mem[912] = -3'h1;
         mem[913] = -3'h1;
         mem[914] = -3'h1;
         mem[915] = -3'h1;
         mem[916] = -3'h1;
         mem[917] = -3'h1;
         mem[918] = -3'h1;
         mem[919] = -3'h1;
         mem[920] = -3'h1;
         mem[921] = -3'h1;
         mem[922] = -3'h1;
         mem[923] = -3'h1;
         mem[924] = -3'h1;
         mem[925] = -3'h1;
         mem[926] = -3'h1;
         mem[927] = -3'h1;
         mem[928] = -3'h1;
         mem[929] = -3'h1;
         mem[930] = -3'h1;
         mem[931] = -3'h1;
         mem[932] = -3'h1;
         mem[933] = -3'h1;
         mem[934] = -3'h1;
         mem[935] = -3'h1;
         mem[936] = -3'h1;
         mem[937] = -3'h1;
         mem[938] = -3'h1;
         mem[939] = -3'h1;
         mem[940] = -3'h1;
         mem[941] = -3'h1;
         mem[942] = -3'h1;
         mem[943] = -3'h1;
         mem[944] = -3'h1;
         mem[945] = -3'h1;
         mem[946] = -3'h1;
         mem[947] = -3'h1;
         mem[948] = -3'h1;
         mem[949] = -3'h1;
         mem[950] = -3'h1;
         mem[951] = -3'h1;
         mem[952] = -3'h1;
         mem[953] = -3'h1;
         mem[954] = -3'h1;
         mem[955] = -3'h1;
         mem[956] = -3'h1;
         mem[957] = -3'h1;
         mem[958] = -3'h1;
         mem[959] = -3'h1;
         mem[960] = -3'h1;
         mem[961] = -3'h1;
         mem[962] = -3'h1;
         mem[963] = -3'h1;
         mem[964] = -3'h1;
         mem[965] = -3'h1;
         mem[966] = -3'h1;
         mem[967] = -3'h1;
         mem[968] = -3'h1;
         mem[969] = -3'h1;
         mem[970] = -3'h1;
         mem[971] = -3'h1;
         mem[972] = -3'h1;
         mem[973] = -3'h1;
         mem[974] = -3'h1;
         mem[975] = -3'h1;
         mem[976] = -3'h1;
         mem[977] = -3'h1;
         mem[978] = -3'h1;
         mem[979] = -3'h1;
         mem[980] = -3'h1;
         mem[981] = -3'h1;
         mem[982] = -3'h1;
         mem[983] = -3'h1;
         mem[984] = -3'h1;
         mem[985] = -3'h1;
         mem[986] = -3'h1;
         mem[987] = -3'h1;
         mem[988] = -3'h1;
         mem[989] = -3'h1;
         mem[990] = -3'h1;
         mem[991] = -3'h1;
         mem[992] = -3'h1;
         mem[993] = -3'h1;
         mem[994] = -3'h1;
         mem[995] = -3'h1;
         mem[996] = -3'h1;
         mem[997] = -3'h1;
         mem[998] = -3'h1;
         mem[999] = -3'h1;
         mem[1000] = -3'h1;
         mem[1001] = -3'h1;
         mem[1002] = -3'h1;
         mem[1003] = -3'h1;
         mem[1004] = -3'h1;
         mem[1005] = -3'h1;
         mem[1006] = -3'h1;
         mem[1007] = -3'h1;
         mem[1008] = -3'h1;
         mem[1009] = -3'h1;
         mem[1010] = -3'h1;
         mem[1011] = -3'h1;
         mem[1012] = -3'h1;
         mem[1013] = -3'h1;
         mem[1014] = -3'h1;
         mem[1015] = -3'h1;
         mem[1016] = -3'h1;
         mem[1017] = -3'h1;
         mem[1018] = -3'h1;
         mem[1019] = -3'h1;
         mem[1020] = -3'h1;
         mem[1021] = -3'h1;
         mem[1022] = -3'h1;
         mem[1023] = -3'h1;
         mem[1024] = -3'h1;
         mem[1025] = -3'h1;
         mem[1026] = -3'h1;
         mem[1027] = -3'h1;
         mem[1028] = -3'h1;
         mem[1029] = -3'h1;
         mem[1030] = -3'h1;
         mem[1031] = -3'h1;
         mem[1032] = -3'h1;
         mem[1033] = -3'h1;
         mem[1034] = -3'h1;
         mem[1035] = -3'h1;
         mem[1036] = -3'h1;
         mem[1037] = -3'h1;
         mem[1038] = -3'h1;
         mem[1039] = -3'h1;
         mem[1040] = -3'h1;
         mem[1041] = -3'h1;
         mem[1042] = -3'h1;
         mem[1043] = -3'h1;
         mem[1044] = -3'h1;
         mem[1045] = -3'h1;
         mem[1046] = -3'h1;
         mem[1047] = -3'h1;
         mem[1048] = -3'h1;
         mem[1049] = -3'h1;
         mem[1050] = -3'h1;
         mem[1051] = -3'h1;
         mem[1052] = -3'h1;
         mem[1053] = -3'h1;
         mem[1054] = -3'h1;
         mem[1055] = -3'h1;
         mem[1056] = -3'h1;
         mem[1057] = -3'h1;
         mem[1058] = -3'h1;
         mem[1059] = -3'h1;
         mem[1060] = -3'h1;
         mem[1061] = -3'h1;
         mem[1062] = -3'h1;
         mem[1063] = -3'h1;
         mem[1064] = -3'h1;
         mem[1065] = -3'h1;
         mem[1066] = -3'h1;
         mem[1067] = -3'h1;
         mem[1068] = -3'h1;
         mem[1069] = -3'h1;
         mem[1070] = -3'h1;
         mem[1071] = -3'h1;
         mem[1072] = -3'h1;
         mem[1073] = -3'h1;
         mem[1074] = -3'h1;
         mem[1075] = -3'h1;
         mem[1076] = -3'h1;
         mem[1077] = -3'h1;
         mem[1078] = -3'h1;
         mem[1079] = -3'h1;
         mem[1080] = -3'h1;
         mem[1081] = -3'h1;
         mem[1082] = -3'h1;
         mem[1083] = -3'h1;
         mem[1084] = -3'h1;
         mem[1085] = -3'h1;
         mem[1086] = -3'h1;
         mem[1087] = -3'h1;
         mem[1088] = -3'h1;
         mem[1089] = -3'h1;
         mem[1090] = -3'h1;
         mem[1091] = -3'h1;
         mem[1092] = -3'h1;
         mem[1093] = -3'h1;
         mem[1094] = -3'h1;
         mem[1095] = -3'h1;
         mem[1096] = -3'h1;
         mem[1097] = -3'h1;
         mem[1098] = -3'h1;
         mem[1099] = -3'h1;
         mem[1100] = -3'h1;
         mem[1101] = -3'h1;
         mem[1102] = -3'h1;
         mem[1103] = -3'h1;
         mem[1104] = -3'h1;
         mem[1105] = -3'h1;
         mem[1106] = -3'h1;
         mem[1107] = -3'h1;
         mem[1108] = -3'h1;
         mem[1109] = -3'h1;
         mem[1110] = -3'h1;
         mem[1111] = -3'h1;
         mem[1112] = -3'h1;
         mem[1113] = -3'h1;
         mem[1114] = -3'h1;
         mem[1115] = -3'h1;
         mem[1116] = -3'h1;
         mem[1117] = -3'h1;
         mem[1118] = -3'h1;
         mem[1119] = -3'h1;
         mem[1120] = -3'h1;
         mem[1121] = -3'h1;
         mem[1122] = -3'h1;
         mem[1123] = -3'h1;
         mem[1124] = -3'h1;
         mem[1125] = -3'h1;
         mem[1126] = -3'h1;
         mem[1127] = -3'h1;
         mem[1128] = -3'h1;
         mem[1129] = -3'h1;
         mem[1130] = -3'h1;
         mem[1131] = -3'h1;
         mem[1132] = -3'h1;
         mem[1133] = -3'h1;
         mem[1134] = -3'h1;
         mem[1135] = -3'h1;
         mem[1136] = -3'h1;
         mem[1137] = -3'h1;
         mem[1138] = -3'h1;
         mem[1139] = -3'h1;
         mem[1140] = -3'h1;
         mem[1141] = -3'h1;
         mem[1142] = -3'h1;
         mem[1143] = -3'h1;
         mem[1144] = -3'h1;
         mem[1145] = -3'h1;
         mem[1146] = -3'h1;
         mem[1147] = -3'h1;
         mem[1148] = -3'h1;
         mem[1149] = -3'h1;
         mem[1150] = -3'h1;
         mem[1151] = -3'h1;
         mem[1152] = -3'h1;
         mem[1153] = -3'h1;
         mem[1154] = -3'h1;
         mem[1155] = -3'h1;
         mem[1156] = -3'h1;
         mem[1157] = -3'h1;
         mem[1158] = -3'h1;
         mem[1159] = -3'h1;
         mem[1160] = -3'h1;
         mem[1161] = -3'h1;
         mem[1162] = -3'h1;
         mem[1163] = -3'h1;
         mem[1164] = -3'h1;
         mem[1165] = -3'h1;
         mem[1166] = -3'h1;
         mem[1167] = -3'h1;
         mem[1168] = -3'h1;
         mem[1169] = -3'h1;
         mem[1170] = -3'h1;
         mem[1171] = -3'h1;
         mem[1172] = -3'h1;
         mem[1173] = -3'h1;
         mem[1174] = -3'h1;
         mem[1175] = -3'h1;
         mem[1176] = -3'h1;
         mem[1177] = -3'h1;
         mem[1178] = -3'h1;
         mem[1179] = -3'h1;
         mem[1180] = -3'h1;
         mem[1181] = -3'h1;
         mem[1182] = -3'h1;
         mem[1183] = -3'h1;
         mem[1184] = -3'h1;
         mem[1185] = -3'h1;
         mem[1186] = -3'h1;
         mem[1187] = -3'h1;
         mem[1188] = -3'h1;
         mem[1189] = -3'h1;
         mem[1190] = -3'h1;
         mem[1191] = -3'h1;
         mem[1192] = -3'h1;
         mem[1193] = -3'h1;
         mem[1194] = -3'h1;
         mem[1195] = -3'h1;
         mem[1196] = -3'h1;
         mem[1197] = -3'h1;
         mem[1198] = -3'h1;
         mem[1199] = -3'h1;
         mem[1200] = -3'h1;
         mem[1201] = -3'h1;
         mem[1202] = -3'h1;
         mem[1203] = -3'h1;
         mem[1204] = -3'h1;
         mem[1205] = -3'h1;
         mem[1206] = -3'h1;
         mem[1207] = -3'h1;
         mem[1208] = -3'h1;
         mem[1209] = -3'h1;
         mem[1210] = -3'h1;
         mem[1211] = -3'h1;
         mem[1212] = -3'h1;
         mem[1213] = -3'h1;
         mem[1214] = -3'h1;
         mem[1215] = -3'h1;
         mem[1216] = -3'h1;
         mem[1217] = -3'h1;
         mem[1218] = -3'h1;
         mem[1219] = -3'h1;
         mem[1220] = -3'h1;
         mem[1221] = -3'h1;
         mem[1222] = -3'h1;
         mem[1223] = -3'h1;
         mem[1224] = -3'h1;
         mem[1225] = -3'h1;
         mem[1226] = -3'h1;
         mem[1227] = -3'h1;
         mem[1228] = -3'h1;
         mem[1229] = -3'h1;
         mem[1230] = -3'h1;
         mem[1231] = -3'h1;
         mem[1232] = -3'h1;
         mem[1233] = -3'h1;
         mem[1234] = -3'h1;
         mem[1235] = -3'h1;
         mem[1236] = -3'h1;
         mem[1237] = -3'h1;
         mem[1238] = -3'h1;
         mem[1239] = -3'h1;
         mem[1240] = -3'h1;
         mem[1241] = -3'h1;
         mem[1242] = -3'h1;
         mem[1243] = -3'h1;
         mem[1244] = -3'h1;
         mem[1245] = -3'h1;
         mem[1246] = -3'h1;
         mem[1247] = -3'h1;
         mem[1248] = -3'h1;
         mem[1249] = -3'h1;
         mem[1250] = -3'h1;
         mem[1251] = -3'h1;
         mem[1252] = -3'h1;
         mem[1253] = -3'h1;
         mem[1254] = -3'h1;
         mem[1255] = -3'h1;
         mem[1256] = -3'h1;
         mem[1257] = -3'h1;
         mem[1258] = -3'h1;
         mem[1259] = -3'h1;
         mem[1260] = -3'h1;
         mem[1261] = -3'h1;
         mem[1262] = -3'h1;
         mem[1263] = -3'h1;
         mem[1264] = -3'h1;
         mem[1265] = -3'h1;
         mem[1266] = -3'h1;
         mem[1267] = -3'h1;
         mem[1268] = -3'h1;
         mem[1269] = -3'h1;
         mem[1270] = -3'h1;
         mem[1271] = -3'h1;
         mem[1272] = -3'h1;
         mem[1273] = -3'h1;
         mem[1274] = -3'h1;
         mem[1275] = -3'h1;
         mem[1276] = -3'h1;
         mem[1277] = -3'h1;
         mem[1278] = -3'h1;
         mem[1279] = -3'h1;
         mem[1280] = -3'h1;
         mem[1281] = -3'h1;
         mem[1282] = -3'h1;
         mem[1283] = -3'h1;
         mem[1284] = -3'h1;
         mem[1285] = -3'h1;
         mem[1286] = -3'h1;
         mem[1287] = -3'h1;
         mem[1288] = -3'h1;
         mem[1289] = -3'h1;
         mem[1290] = -3'h1;
         mem[1291] = -3'h1;
         mem[1292] = -3'h1;
         mem[1293] = -3'h1;
         mem[1294] = -3'h1;
         mem[1295] = -3'h1;
         mem[1296] = -3'h1;
         mem[1297] = -3'h1;
         mem[1298] = -3'h1;
         mem[1299] = -3'h1;
         mem[1300] = -3'h1;
         mem[1301] = -3'h1;
         mem[1302] = -3'h1;
         mem[1303] = -3'h1;
         mem[1304] = -3'h1;
         mem[1305] = -3'h1;
         mem[1306] = -3'h1;
         mem[1307] = -3'h1;
         mem[1308] = -3'h1;
         mem[1309] = -3'h1;
         mem[1310] = -3'h1;
         mem[1311] = -3'h1;
         mem[1312] = -3'h1;
         mem[1313] = -3'h1;
         mem[1314] = -3'h1;
         mem[1315] = -3'h1;
         mem[1316] = -3'h1;
         mem[1317] = -3'h1;
         mem[1318] = -3'h1;
         mem[1319] = -3'h1;
         mem[1320] = -3'h1;
         mem[1321] = -3'h1;
         mem[1322] = -3'h1;
         mem[1323] = -3'h1;
         mem[1324] = -3'h1;
         mem[1325] = -3'h1;
         mem[1326] = -3'h1;
         mem[1327] = -3'h1;
         mem[1328] = -3'h1;
         mem[1329] = -3'h1;
         mem[1330] = -3'h1;
         mem[1331] = -3'h1;
         mem[1332] = -3'h1;
         mem[1333] = -3'h1;
         mem[1334] = -3'h1;
         mem[1335] = -3'h1;
         mem[1336] = -3'h1;
         mem[1337] = -3'h1;
         mem[1338] = -3'h1;
         mem[1339] = -3'h1;
         mem[1340] = -3'h1;
         mem[1341] = -3'h1;
         mem[1342] = -3'h1;
         mem[1343] = -3'h1;
         mem[1344] = -3'h1;
         mem[1345] = -3'h1;
         mem[1346] = -3'h1;
         mem[1347] = -3'h1;
         mem[1348] = -3'h1;
         mem[1349] = -3'h1;
         mem[1350] = -3'h1;
         mem[1351] = -3'h1;
         mem[1352] = -3'h1;
         mem[1353] = -3'h1;
         mem[1354] = -3'h1;
         mem[1355] = -3'h1;
         mem[1356] = -3'h1;
         mem[1357] = -3'h1;
         mem[1358] = -3'h1;
         mem[1359] = -3'h1;
         mem[1360] = -3'h1;
         mem[1361] = -3'h1;
         mem[1362] = -3'h1;
         mem[1363] = -3'h1;
         mem[1364] = -3'h1;
         mem[1365] = -3'h1;
         mem[1366] = -3'h1;
         mem[1367] = -3'h1;
         mem[1368] = -3'h1;
         mem[1369] = -3'h1;
         mem[1370] = -3'h1;
         mem[1371] = -3'h1;
         mem[1372] = -3'h1;
         mem[1373] = -3'h1;
         mem[1374] = -3'h1;
         mem[1375] = -3'h1;
         mem[1376] = -3'h1;
         mem[1377] = -3'h1;
         mem[1378] = -3'h1;
         mem[1379] = -3'h1;
         mem[1380] = -3'h1;
         mem[1381] = -3'h1;
         mem[1382] = -3'h1;
         mem[1383] = -3'h1;
         mem[1384] = -3'h1;
         mem[1385] = -3'h1;
         mem[1386] = -3'h1;
         mem[1387] = -3'h1;
         mem[1388] = -3'h1;
         mem[1389] = -3'h1;
         mem[1390] = -3'h1;
         mem[1391] = -3'h1;
         mem[1392] = -3'h1;
         mem[1393] = -3'h1;
         mem[1394] = -3'h1;
         mem[1395] = -3'h1;
         mem[1396] = -3'h1;
         mem[1397] = -3'h1;
         mem[1398] = -3'h1;
         mem[1399] = -3'h1;
         mem[1400] = -3'h1;
         mem[1401] = -3'h1;
         mem[1402] = -3'h1;
         mem[1403] = -3'h1;
         mem[1404] = -3'h1;
         mem[1405] = -3'h1;
         mem[1406] = -3'h1;
         mem[1407] = -3'h1;
         mem[1408] = -3'h1;
         mem[1409] = -3'h1;
         mem[1410] = -3'h1;
         mem[1411] = -3'h1;
         mem[1412] = -3'h1;
         mem[1413] = -3'h1;
         mem[1414] = -3'h1;
         mem[1415] = -3'h1;
         mem[1416] = -3'h1;
         mem[1417] = -3'h1;
         mem[1418] = -3'h1;
         mem[1419] = -3'h1;
         mem[1420] = -3'h1;
         mem[1421] = -3'h1;
         mem[1422] = -3'h1;
         mem[1423] = -3'h1;
         mem[1424] = -3'h1;
         mem[1425] = -3'h1;
         mem[1426] = -3'h1;
         mem[1427] = -3'h1;
         mem[1428] = -3'h1;
         mem[1429] = -3'h1;
         mem[1430] = -3'h1;
         mem[1431] = -3'h1;
         mem[1432] = -3'h1;
         mem[1433] = -3'h1;
         mem[1434] = -3'h1;
         mem[1435] = -3'h1;
         mem[1436] = -3'h1;
         mem[1437] = -3'h1;
         mem[1438] = -3'h1;
         mem[1439] = -3'h1;
         mem[1440] = -3'h1;
         mem[1441] = -3'h1;
         mem[1442] = -3'h1;
         mem[1443] = -3'h1;
         mem[1444] = -3'h1;
         mem[1445] = -3'h1;
         mem[1446] = -3'h1;
         mem[1447] = -3'h1;
         mem[1448] = -3'h1;
         mem[1449] = -3'h1;
         mem[1450] = -3'h1;
         mem[1451] = -3'h1;
         mem[1452] = -3'h1;
         mem[1453] = -3'h1;
         mem[1454] = -3'h1;
         mem[1455] = -3'h1;
         mem[1456] = -3'h1;
         mem[1457] = -3'h1;
         mem[1458] = -3'h1;
         mem[1459] = -3'h1;
         mem[1460] = -3'h1;
         mem[1461] = -3'h1;
         mem[1462] = -3'h1;
         mem[1463] = -3'h1;
         mem[1464] = -3'h1;
         mem[1465] = -3'h1;
         mem[1466] = -3'h1;
         mem[1467] = -3'h1;
         mem[1468] = -3'h1;
         mem[1469] = -3'h1;
         mem[1470] = -3'h1;
         mem[1471] = -3'h1;
         mem[1472] = -3'h1;
         mem[1473] = -3'h1;
         mem[1474] = -3'h1;
         mem[1475] = -3'h1;
         mem[1476] = -3'h1;
         mem[1477] = -3'h1;
         mem[1478] = -3'h1;
         mem[1479] = -3'h1;
         mem[1480] = -3'h1;
         mem[1481] = -3'h1;
         mem[1482] = -3'h1;
         mem[1483] = -3'h1;
         mem[1484] = -3'h1;
         mem[1485] = -3'h1;
         mem[1486] = -3'h1;
         mem[1487] = -3'h1;
         mem[1488] = -3'h1;
         mem[1489] = -3'h1;
         mem[1490] = -3'h1;
         mem[1491] = -3'h1;
         mem[1492] = -3'h1;
         mem[1493] = -3'h1;
         mem[1494] = -3'h1;
         mem[1495] = -3'h1;
         mem[1496] = -3'h1;
         mem[1497] = -3'h1;
         mem[1498] = -3'h1;
         mem[1499] = -3'h1;
         mem[1500] = -3'h1;
         mem[1501] = -3'h1;
         mem[1502] = -3'h1;
         mem[1503] = -3'h1;
         mem[1504] = -3'h1;
         mem[1505] = -3'h1;
         mem[1506] = -3'h1;
         mem[1507] = -3'h1;
         mem[1508] = -3'h1;
         mem[1509] = -3'h1;
         mem[1510] = -3'h1;
         mem[1511] = -3'h1;
         mem[1512] = -3'h1;
         mem[1513] = -3'h1;
         mem[1514] = -3'h1;
         mem[1515] = -3'h1;
         mem[1516] = -3'h1;
         mem[1517] = -3'h1;
         mem[1518] = -3'h1;
         mem[1519] = -3'h1;
         mem[1520] = -3'h1;
         mem[1521] = -3'h1;
         mem[1522] = -3'h1;
         mem[1523] = -3'h1;
         mem[1524] = -3'h1;
         mem[1525] = -3'h1;
         mem[1526] = -3'h1;
         mem[1527] = -3'h1;
         mem[1528] = -3'h1;
         mem[1529] = -3'h1;
         mem[1530] = -3'h1;
         mem[1531] = -3'h1;
         mem[1532] = -3'h1;
         mem[1533] = -3'h1;
         mem[1534] = -3'h1;
         mem[1535] = -3'h1;
         mem[1536] = -3'h1;
         mem[1537] = -3'h1;
         mem[1538] = -3'h1;
         mem[1539] = -3'h1;
         mem[1540] = -3'h1;
         mem[1541] = -3'h1;
         mem[1542] = -3'h1;
         mem[1543] = -3'h1;
         mem[1544] = -3'h1;
         mem[1545] = -3'h1;
         mem[1546] = -3'h1;
         mem[1547] = -3'h1;
         mem[1548] = -3'h1;
         mem[1549] = -3'h1;
         mem[1550] = -3'h1;
         mem[1551] = -3'h1;
         mem[1552] = -3'h1;
         mem[1553] = -3'h1;
         mem[1554] = -3'h1;
         mem[1555] = -3'h1;
         mem[1556] = -3'h1;
         mem[1557] = -3'h1;
         mem[1558] = -3'h1;
         mem[1559] = -3'h1;
         mem[1560] = -3'h1;
         mem[1561] = -3'h1;
         mem[1562] = -3'h1;
         mem[1563] = -3'h1;
         mem[1564] = -3'h1;
         mem[1565] = -3'h1;
         mem[1566] = -3'h1;
         mem[1567] = -3'h1;
         mem[1568] = -3'h1;
         mem[1569] = -3'h1;
         mem[1570] = -3'h1;
         mem[1571] = -3'h1;
         mem[1572] = -3'h1;
         mem[1573] = -3'h1;
         mem[1574] = -3'h1;
         mem[1575] = -3'h1;
         mem[1576] = -3'h1;
         mem[1577] = -3'h1;
         mem[1578] = -3'h1;
         mem[1579] = -3'h1;
         mem[1580] = -3'h1;
         mem[1581] = -3'h1;
         mem[1582] = -3'h1;
         mem[1583] = -3'h1;
         mem[1584] = -3'h1;
         mem[1585] = -3'h1;
         mem[1586] = -3'h1;
         mem[1587] = -3'h1;
         mem[1588] = -3'h1;
         mem[1589] = -3'h1;
         mem[1590] = -3'h1;
         mem[1591] = -3'h1;
         mem[1592] = -3'h1;
         mem[1593] = -3'h1;
         mem[1594] = -3'h1;
         mem[1595] = -3'h1;
         mem[1596] = -3'h1;
         mem[1597] = -3'h1;
         mem[1598] = -3'h1;
         mem[1599] = -3'h1;
         mem[1600] = -3'h1;
         mem[1601] = -3'h1;
         mem[1602] = -3'h1;
         mem[1603] = -3'h1;
         mem[1604] = -3'h1;
         mem[1605] = -3'h1;
         mem[1606] = -3'h1;
         mem[1607] = -3'h1;
         mem[1608] = -3'h1;
         mem[1609] = -3'h1;
         mem[1610] = -3'h1;
         mem[1611] = -3'h1;
         mem[1612] = -3'h1;
         mem[1613] = -3'h1;
         mem[1614] = -3'h1;
         mem[1615] = -3'h1;
         mem[1616] = -3'h1;
         mem[1617] = -3'h1;
         mem[1618] = -3'h1;
         mem[1619] = -3'h1;
         mem[1620] = -3'h1;
         mem[1621] = -3'h1;
         mem[1622] = -3'h1;
         mem[1623] = -3'h1;
         mem[1624] = -3'h1;
         mem[1625] = -3'h1;
         mem[1626] = -3'h1;
         mem[1627] = -3'h1;
         mem[1628] = -3'h1;
         mem[1629] = -3'h1;
         mem[1630] = -3'h1;
         mem[1631] = -3'h1;
         mem[1632] = -3'h1;
         mem[1633] = -3'h1;
         mem[1634] = -3'h1;
         mem[1635] = -3'h1;
         mem[1636] = -3'h1;
         mem[1637] = -3'h1;
         mem[1638] = -3'h1;
         mem[1639] = -3'h1;
         mem[1640] = -3'h1;
         mem[1641] = -3'h1;
         mem[1642] = -3'h1;
         mem[1643] = -3'h1;
         mem[1644] = -3'h1;
         mem[1645] = -3'h1;
         mem[1646] = -3'h1;
         mem[1647] = -3'h1;
         mem[1648] = -3'h1;
         mem[1649] = -3'h1;
         mem[1650] = -3'h1;
         mem[1651] = -3'h1;
         mem[1652] = -3'h1;
         mem[1653] = -3'h1;
         mem[1654] = -3'h1;
         mem[1655] = -3'h1;
         mem[1656] = -3'h1;
         mem[1657] = -3'h1;
         mem[1658] = -3'h1;
         mem[1659] = -3'h1;
         mem[1660] = -3'h1;
         mem[1661] = -3'h1;
         mem[1662] = -3'h1;
         mem[1663] = -3'h1;
         mem[1664] = -3'h1;
         mem[1665] = -3'h1;
         mem[1666] = -3'h1;
         mem[1667] = -3'h1;
         mem[1668] = -3'h1;
         mem[1669] = -3'h1;
         mem[1670] = -3'h1;
         mem[1671] = -3'h1;
         mem[1672] = -3'h1;
         mem[1673] = -3'h1;
         mem[1674] = -3'h1;
         mem[1675] = -3'h1;
         mem[1676] = -3'h1;
         mem[1677] = -3'h1;
         mem[1678] = -3'h1;
         mem[1679] = -3'h1;
         mem[1680] = -3'h1;
         mem[1681] = -3'h1;
         mem[1682] = -3'h1;
         mem[1683] = -3'h1;
         mem[1684] = -3'h1;
         mem[1685] = -3'h1;
         mem[1686] = -3'h1;
         mem[1687] = -3'h1;
         mem[1688] = -3'h1;
         mem[1689] = -3'h1;
         mem[1690] = -3'h1;
         mem[1691] = -3'h1;
         mem[1692] = -3'h1;
         mem[1693] = -3'h1;
         mem[1694] = -3'h1;
         mem[1695] = -3'h1;
         mem[1696] = -3'h1;
         mem[1697] = -3'h1;
         mem[1698] = -3'h1;
         mem[1699] = -3'h1;
         mem[1700] = -3'h1;
         mem[1701] = -3'h1;
         mem[1702] = -3'h1;
         mem[1703] = -3'h1;
         mem[1704] = -3'h1;
         mem[1705] = -3'h1;
         mem[1706] = -3'h1;
         mem[1707] = -3'h1;
         mem[1708] = -3'h1;
         mem[1709] = -3'h1;
         mem[1710] = -3'h1;
         mem[1711] = -3'h1;
         mem[1712] = -3'h1;
         mem[1713] = -3'h1;
         mem[1714] = -3'h1;
         mem[1715] = -3'h1;
         mem[1716] = -3'h1;
         mem[1717] = -3'h1;
         mem[1718] = -3'h1;
         mem[1719] = -3'h1;
         mem[1720] = -3'h1;
         mem[1721] = -3'h1;
         mem[1722] = -3'h1;
         mem[1723] = -3'h1;
         mem[1724] = -3'h1;
         mem[1725] = -3'h1;
         mem[1726] = -3'h1;
         mem[1727] = -3'h1;
         mem[1728] = -3'h1;
         mem[1729] = -3'h1;
         mem[1730] = -3'h1;
         mem[1731] = -3'h1;
         mem[1732] = -3'h1;
         mem[1733] = -3'h1;
         mem[1734] = -3'h1;
         mem[1735] = -3'h1;
         mem[1736] = -3'h1;
         mem[1737] = -3'h1;
         mem[1738] = -3'h1;
         mem[1739] = -3'h1;
         mem[1740] = -3'h1;
         mem[1741] = -3'h1;
         mem[1742] = -3'h1;
         mem[1743] = -3'h1;
         mem[1744] = -3'h1;
         mem[1745] = -3'h1;
         mem[1746] = -3'h1;
         mem[1747] = -3'h1;
         mem[1748] = -3'h1;
         mem[1749] = -3'h1;
         mem[1750] = -3'h1;
         mem[1751] = -3'h1;
         mem[1752] = -3'h1;
         mem[1753] = -3'h1;
         mem[1754] = -3'h1;
         mem[1755] = -3'h1;
         mem[1756] = -3'h1;
         mem[1757] = -3'h1;
         mem[1758] = -3'h1;
         mem[1759] = -3'h1;
         mem[1760] = -3'h1;
         mem[1761] = -3'h1;
         mem[1762] = -3'h1;
         mem[1763] = -3'h1;
         mem[1764] = -3'h1;
         mem[1765] = -3'h1;
         mem[1766] = -3'h1;
         mem[1767] = -3'h1;
         mem[1768] = -3'h1;
         mem[1769] = -3'h1;
         mem[1770] = -3'h1;
         mem[1771] = -3'h1;
         mem[1772] = -3'h1;
         mem[1773] = -3'h1;
         mem[1774] = -3'h1;
         mem[1775] = -3'h1;
         mem[1776] = -3'h1;
         mem[1777] = -3'h1;
         mem[1778] = -3'h1;
         mem[1779] = -3'h1;
         mem[1780] = -3'h1;
         mem[1781] = -3'h1;
         mem[1782] = -3'h1;
         mem[1783] = -3'h1;
         mem[1784] = -3'h1;
         mem[1785] = -3'h1;
         mem[1786] = -3'h1;
         mem[1787] = -3'h1;
         mem[1788] = -3'h1;
         mem[1789] = -3'h1;
         mem[1790] = -3'h1;
         mem[1791] = -3'h1;
         mem[1792] = -3'h1;
         mem[1793] = -3'h1;
         mem[1794] = -3'h1;
         mem[1795] = -3'h1;
         mem[1796] = -3'h1;
         mem[1797] = -3'h1;
         mem[1798] = -3'h1;
         mem[1799] = -3'h1;
         mem[1800] = -3'h1;
         mem[1801] = -3'h1;
         mem[1802] = -3'h1;
         mem[1803] = -3'h1;
         mem[1804] = -3'h1;
         mem[1805] = -3'h1;
         mem[1806] = -3'h1;
         mem[1807] = -3'h1;
         mem[1808] = -3'h1;
         mem[1809] = -3'h1;
         mem[1810] = -3'h1;
         mem[1811] = -3'h1;
         mem[1812] = -3'h1;
         mem[1813] = -3'h1;
         mem[1814] = -3'h1;
         mem[1815] = -3'h1;
         mem[1816] = -3'h1;
         mem[1817] = -3'h1;
         mem[1818] = -3'h1;
         mem[1819] = -3'h1;
         mem[1820] = -3'h1;
         mem[1821] = -3'h1;
         mem[1822] = -3'h1;
         mem[1823] = -3'h1;
         mem[1824] = -3'h1;
         mem[1825] = -3'h1;
         mem[1826] = -3'h1;
         mem[1827] = -3'h1;
         mem[1828] = -3'h1;
         mem[1829] = -3'h1;
         mem[1830] = -3'h1;
         mem[1831] = -3'h1;
         mem[1832] = -3'h1;
         mem[1833] = -3'h1;
         mem[1834] = -3'h1;
         mem[1835] = -3'h1;
         mem[1836] = -3'h1;
         mem[1837] = -3'h1;
         mem[1838] = -3'h1;
         mem[1839] = -3'h1;
         mem[1840] = -3'h1;
         mem[1841] = -3'h1;
         mem[1842] = -3'h1;
         mem[1843] = -3'h1;
         mem[1844] = -3'h1;
         mem[1845] = -3'h1;
         mem[1846] = -3'h1;
         mem[1847] = -3'h1;
         mem[1848] = -3'h1;
         mem[1849] = -3'h1;
         mem[1850] = -3'h1;
         mem[1851] = -3'h1;
         mem[1852] = -3'h1;
         mem[1853] = -3'h1;
         mem[1854] = -3'h1;
         mem[1855] = -3'h1;
         mem[1856] = -3'h1;
         mem[1857] = -3'h1;
         mem[1858] = -3'h1;
         mem[1859] = -3'h1;
         mem[1860] = -3'h1;
         mem[1861] = -3'h1;
         mem[1862] = -3'h1;
         mem[1863] = -3'h1;
         mem[1864] = -3'h1;
         mem[1865] = -3'h1;
         mem[1866] = -3'h1;
         mem[1867] = -3'h1;
         mem[1868] = -3'h1;
         mem[1869] = -3'h1;
         mem[1870] = -3'h1;
         mem[1871] = -3'h1;
         mem[1872] = -3'h1;
         mem[1873] = -3'h1;
         mem[1874] = -3'h1;
         mem[1875] = -3'h1;
         mem[1876] = -3'h1;
         mem[1877] = -3'h1;
         mem[1878] = -3'h1;
         mem[1879] = -3'h1;
         mem[1880] = -3'h1;
         mem[1881] = -3'h1;
         mem[1882] = -3'h1;
         mem[1883] = -3'h1;
         mem[1884] = -3'h1;
         mem[1885] = -3'h1;
         mem[1886] = -3'h1;
         mem[1887] = -3'h1;
         mem[1888] = -3'h1;
         mem[1889] = -3'h1;
         mem[1890] = -3'h1;
         mem[1891] = -3'h1;
         mem[1892] = -3'h1;
         mem[1893] = -3'h1;
         mem[1894] = -3'h1;
         mem[1895] = -3'h1;
         mem[1896] = -3'h1;
         mem[1897] = -3'h1;
         mem[1898] = -3'h1;
         mem[1899] = -3'h1;
         mem[1900] = -3'h1;
         mem[1901] = -3'h1;
         mem[1902] = -3'h1;
         mem[1903] = -3'h1;
         mem[1904] = -3'h1;
         mem[1905] = -3'h1;
         mem[1906] = -3'h1;
         mem[1907] = -3'h1;
         mem[1908] = -3'h1;
         mem[1909] = -3'h1;
         mem[1910] = -3'h1;
         mem[1911] = -3'h1;
         mem[1912] = -3'h1;
         mem[1913] = -3'h1;
         mem[1914] = -3'h1;
         mem[1915] = -3'h1;
         mem[1916] = -3'h1;
         mem[1917] = -3'h1;
         mem[1918] = -3'h1;
         mem[1919] = -3'h1;
         mem[1920] = -3'h1;
         mem[1921] = -3'h1;
         mem[1922] = -3'h1;
         mem[1923] = -3'h1;
         mem[1924] = -3'h1;
         mem[1925] = -3'h1;
         mem[1926] = -3'h1;
         mem[1927] = -3'h1;
         mem[1928] = -3'h1;
         mem[1929] = -3'h1;
         mem[1930] = -3'h1;
         mem[1931] = -3'h1;
         mem[1932] = -3'h1;
         mem[1933] = -3'h1;
         mem[1934] = -3'h1;
         mem[1935] = -3'h1;
         mem[1936] = -3'h1;
         mem[1937] = -3'h1;
         mem[1938] = -3'h1;
         mem[1939] = -3'h1;
         mem[1940] = -3'h1;
         mem[1941] = -3'h1;
         mem[1942] = -3'h1;
         mem[1943] = -3'h1;
         mem[1944] = -3'h1;
         mem[1945] = -3'h1;
         mem[1946] = -3'h1;
         mem[1947] = -3'h1;
         mem[1948] = -3'h1;
         mem[1949] = -3'h1;
         mem[1950] = -3'h1;
         mem[1951] = -3'h1;
         mem[1952] = -3'h1;
         mem[1953] = -3'h1;
         mem[1954] = -3'h1;
         mem[1955] = -3'h1;
         mem[1956] = -3'h1;
         mem[1957] = -3'h1;
         mem[1958] = -3'h1;
         mem[1959] = -3'h1;
         mem[1960] = -3'h1;
         mem[1961] = -3'h1;
         mem[1962] = -3'h1;
         mem[1963] = -3'h1;
         mem[1964] = -3'h1;
         mem[1965] = -3'h1;
         mem[1966] = -3'h1;
         mem[1967] = -3'h1;
         mem[1968] = -3'h1;
         mem[1969] = -3'h1;
         mem[1970] = -3'h1;
         mem[1971] = -3'h1;
         mem[1972] = -3'h1;
         mem[1973] = -3'h1;
         mem[1974] = -3'h1;
         mem[1975] = -3'h1;
         mem[1976] = -3'h1;
         mem[1977] = -3'h1;
         mem[1978] = -3'h1;
         mem[1979] = -3'h1;
         mem[1980] = -3'h1;
         mem[1981] = -3'h1;
         mem[1982] = -3'h1;
         mem[1983] = -3'h1;
         mem[1984] = -3'h1;
         mem[1985] = -3'h1;
         mem[1986] = -3'h1;
         mem[1987] = -3'h1;
         mem[1988] = -3'h1;
         mem[1989] = -3'h1;
         mem[1990] = -3'h1;
         mem[1991] = -3'h1;
         mem[1992] = -3'h1;
         mem[1993] = -3'h1;
         mem[1994] = -3'h1;
         mem[1995] = -3'h1;
         mem[1996] = -3'h1;
         mem[1997] = -3'h1;
         mem[1998] = -3'h1;
         mem[1999] = -3'h1;
         mem[2000] = -3'h1;
         mem[2001] = -3'h1;
         mem[2002] = -3'h1;
         mem[2003] = -3'h1;
         mem[2004] = -3'h1;
         mem[2005] = -3'h1;
         mem[2006] = -3'h1;
         mem[2007] = -3'h1;
         mem[2008] = -3'h1;
         mem[2009] = -3'h1;
         mem[2010] = -3'h1;
         mem[2011] = -3'h1;
         mem[2012] = -3'h1;
         mem[2013] = -3'h1;
         mem[2014] = -3'h1;
         mem[2015] = -3'h1;
         mem[2016] = -3'h1;
         mem[2017] = -3'h1;
         mem[2018] = -3'h1;
         mem[2019] = -3'h1;
         mem[2020] = -3'h1;
         mem[2021] = -3'h1;
         mem[2022] = -3'h1;
         mem[2023] = -3'h1;
         mem[2024] = -3'h1;
         mem[2025] = -3'h1;
         mem[2026] = -3'h1;
         mem[2027] = -3'h1;
         mem[2028] = -3'h1;
         mem[2029] = -3'h1;
         mem[2030] = -3'h1;
         mem[2031] = -3'h1;
         mem[2032] = -3'h1;
         mem[2033] = -3'h1;
         mem[2034] = -3'h1;
         mem[2035] = -3'h1;
         mem[2036] = -3'h1;
         mem[2037] = -3'h1;
         mem[2038] = -3'h1;
         mem[2039] = -3'h1;
         mem[2040] = -3'h1;
         mem[2041] = -3'h1;
         mem[2042] = -3'h1;
         mem[2043] = -3'h1;
         mem[2044] = -3'h1;
         mem[2045] = -3'h1;
         mem[2046] = -3'h1;
         mem[2047] = -3'h1;
         mem[2048] = -3'h1;
         mem[2049] = -3'h1;
         mem[2050] = -3'h1;
         mem[2051] = -3'h1;
         mem[2052] = -3'h1;
         mem[2053] = -3'h1;
         mem[2054] = -3'h1;
         mem[2055] = -3'h1;
         mem[2056] = -3'h1;
         mem[2057] = -3'h1;
         mem[2058] = -3'h1;
         mem[2059] = -3'h1;
         mem[2060] = -3'h1;
         mem[2061] = -3'h1;
         mem[2062] = -3'h1;
         mem[2063] = -3'h1;
         mem[2064] = -3'h1;
         mem[2065] = -3'h1;
         mem[2066] = -3'h1;
         mem[2067] = -3'h1;
         mem[2068] = -3'h1;
         mem[2069] = -3'h1;
         mem[2070] = -3'h1;
         mem[2071] = -3'h1;
         mem[2072] = -3'h1;
         mem[2073] = -3'h1;
         mem[2074] = -3'h1;
         mem[2075] = -3'h1;
         mem[2076] = -3'h1;
         mem[2077] = -3'h1;
         mem[2078] = -3'h1;
         mem[2079] = -3'h1;
         mem[2080] = -3'h1;
         mem[2081] = -3'h1;
         mem[2082] = -3'h1;
         mem[2083] = -3'h1;
         mem[2084] = -3'h1;
         mem[2085] = -3'h1;
         mem[2086] = -3'h1;
         mem[2087] = -3'h1;
         mem[2088] = -3'h1;
         mem[2089] = -3'h1;
         mem[2090] = -3'h1;
         mem[2091] = -3'h1;
         mem[2092] = -3'h1;
         mem[2093] = -3'h1;
         mem[2094] = -3'h1;
         mem[2095] = -3'h1;
         mem[2096] = -3'h1;
         mem[2097] = -3'h1;
         mem[2098] = -3'h1;
         mem[2099] = -3'h1;
         mem[2100] = -3'h1;
         mem[2101] = -3'h1;
         mem[2102] = -3'h1;
         mem[2103] = -3'h1;
         mem[2104] = -3'h1;
         mem[2105] = -3'h1;
         mem[2106] = -3'h1;
         mem[2107] = -3'h1;
         mem[2108] = -3'h1;
         mem[2109] = -3'h1;
         mem[2110] = -3'h1;
         mem[2111] = -3'h1;
         mem[2112] = -3'h1;
         mem[2113] = -3'h1;
         mem[2114] = -3'h1;
         mem[2115] = -3'h1;
         mem[2116] = -3'h1;
         mem[2117] = -3'h1;
         mem[2118] = -3'h1;
         mem[2119] = -3'h1;
         mem[2120] = -3'h1;
         mem[2121] = -3'h1;
         mem[2122] = -3'h1;
         mem[2123] = -3'h1;
         mem[2124] = -3'h1;
         mem[2125] = -3'h1;
         mem[2126] = -3'h1;
         mem[2127] = -3'h1;
         mem[2128] = -3'h1;
         mem[2129] = -3'h1;
         mem[2130] = -3'h1;
         mem[2131] = -3'h1;
         mem[2132] = -3'h1;
         mem[2133] = -3'h1;
         mem[2134] = -3'h1;
         mem[2135] = -3'h1;
         mem[2136] = -3'h1;
         mem[2137] = -3'h1;
         mem[2138] = -3'h1;
         mem[2139] = -3'h1;
         mem[2140] = -3'h1;
         mem[2141] = -3'h1;
         mem[2142] = -3'h1;
         mem[2143] = -3'h1;
         mem[2144] = -3'h1;
         mem[2145] = -3'h1;
         mem[2146] = -3'h1;
         mem[2147] = -3'h1;
         mem[2148] = -3'h1;
         mem[2149] = -3'h1;
         mem[2150] = -3'h1;
         mem[2151] = -3'h1;
         mem[2152] = -3'h1;
         mem[2153] = -3'h1;
         mem[2154] = -3'h1;
         mem[2155] = -3'h1;
         mem[2156] = -3'h1;
         mem[2157] = -3'h1;
         mem[2158] = -3'h1;
         mem[2159] = -3'h1;
         mem[2160] = -3'h1;
         mem[2161] = -3'h1;
         mem[2162] = -3'h1;
         mem[2163] = -3'h1;
         mem[2164] = -3'h1;
         mem[2165] = -3'h1;
         mem[2166] = -3'h1;
         mem[2167] = -3'h1;
         mem[2168] = -3'h1;
         mem[2169] = -3'h1;
         mem[2170] = -3'h1;
         mem[2171] = -3'h1;
         mem[2172] = -3'h1;
         mem[2173] = -3'h1;
         mem[2174] = -3'h1;
         mem[2175] = -3'h1;
         mem[2176] = -3'h1;
         mem[2177] = -3'h1;
         mem[2178] = -3'h1;
         mem[2179] = -3'h1;
         mem[2180] = -3'h1;
         mem[2181] = -3'h1;
         mem[2182] = -3'h1;
         mem[2183] = -3'h1;
         mem[2184] = -3'h1;
         mem[2185] = -3'h1;
         mem[2186] = -3'h1;
         mem[2187] = -3'h1;
         mem[2188] = -3'h1;
         mem[2189] = -3'h1;
         mem[2190] = -3'h1;
         mem[2191] = -3'h1;
         mem[2192] = -3'h1;
         mem[2193] = -3'h1;
         mem[2194] = -3'h1;
         mem[2195] = -3'h1;
         mem[2196] = -3'h1;
         mem[2197] = -3'h1;
         mem[2198] = -3'h1;
         mem[2199] = -3'h1;
         mem[2200] = -3'h1;
         mem[2201] = -3'h1;
         mem[2202] = -3'h1;
         mem[2203] = -3'h1;
         mem[2204] = -3'h1;
         mem[2205] = -3'h1;
         mem[2206] = -3'h1;
         mem[2207] = -3'h1;
         mem[2208] = -3'h1;
         mem[2209] = -3'h1;
         mem[2210] = -3'h1;
         mem[2211] = -3'h1;
         mem[2212] = -3'h1;
         mem[2213] = -3'h1;
         mem[2214] = -3'h1;
         mem[2215] = -3'h1;
         mem[2216] = -3'h1;
         mem[2217] = -3'h1;
         mem[2218] = -3'h1;
         mem[2219] = -3'h1;
         mem[2220] = -3'h1;
         mem[2221] = -3'h1;
         mem[2222] = -3'h1;
         mem[2223] = -3'h1;
         mem[2224] = -3'h1;
         mem[2225] = -3'h1;
         mem[2226] = -3'h1;
         mem[2227] = -3'h1;
         mem[2228] = -3'h1;
         mem[2229] = -3'h1;
         mem[2230] = -3'h1;
         mem[2231] = -3'h1;
         mem[2232] = -3'h1;
         mem[2233] = -3'h1;
         mem[2234] = -3'h1;
         mem[2235] = -3'h1;
         mem[2236] = -3'h1;
         mem[2237] = -3'h1;
         mem[2238] = -3'h1;
         mem[2239] = -3'h1;
         mem[2240] = -3'h1;
         mem[2241] = -3'h1;
         mem[2242] = -3'h1;
         mem[2243] = -3'h1;
         mem[2244] = -3'h1;
         mem[2245] = -3'h1;
         mem[2246] = -3'h1;
         mem[2247] = -3'h1;
         mem[2248] = -3'h1;
         mem[2249] = -3'h1;
         mem[2250] = -3'h1;
         mem[2251] = -3'h1;
         mem[2252] = -3'h1;
         mem[2253] = -3'h1;
         mem[2254] = -3'h1;
         mem[2255] = -3'h1;
         mem[2256] = -3'h1;
         mem[2257] = -3'h1;
         mem[2258] = -3'h1;
         mem[2259] = -3'h1;
         mem[2260] = -3'h1;
         mem[2261] = -3'h1;
         mem[2262] = -3'h1;
         mem[2263] = -3'h1;
         mem[2264] = -3'h1;
         mem[2265] = -3'h1;
         mem[2266] = -3'h1;
         mem[2267] = -3'h1;
         mem[2268] = -3'h1;
         mem[2269] = -3'h1;
         mem[2270] = -3'h1;
         mem[2271] = -3'h1;
         mem[2272] = -3'h1;
         mem[2273] = -3'h1;
         mem[2274] = -3'h1;
         mem[2275] = -3'h1;
         mem[2276] = -3'h1;
         mem[2277] = -3'h1;
         mem[2278] = -3'h1;
         mem[2279] = -3'h1;
         mem[2280] = -3'h1;
         mem[2281] = -3'h1;
         mem[2282] = -3'h1;
         mem[2283] = -3'h1;
         mem[2284] = -3'h1;
         mem[2285] = -3'h1;
         mem[2286] = -3'h1;
         mem[2287] = -3'h1;
         mem[2288] = -3'h1;
         mem[2289] = -3'h1;
         mem[2290] = -3'h1;
         mem[2291] = -3'h1;
         mem[2292] = -3'h1;
         mem[2293] = -3'h1;
         mem[2294] = -3'h1;
         mem[2295] = -3'h1;
         mem[2296] = -3'h1;
         mem[2297] = -3'h1;
         mem[2298] = -3'h1;
         mem[2299] = -3'h1;
         mem[2300] = -3'h1;
         mem[2301] = -3'h1;
         mem[2302] = -3'h1;
         mem[2303] = -3'h1;
         mem[2304] = -3'h1;
         mem[2305] = -3'h1;
         mem[2306] = -3'h1;
         mem[2307] = -3'h1;
         mem[2308] = -3'h1;
         mem[2309] = -3'h1;
         mem[2310] = -3'h1;
         mem[2311] = -3'h1;
         mem[2312] = -3'h1;
         mem[2313] = -3'h1;
         mem[2314] = -3'h1;
         mem[2315] = -3'h1;
         mem[2316] = -3'h1;
         mem[2317] = -3'h1;
         mem[2318] = -3'h1;
         mem[2319] = -3'h1;
         mem[2320] = -3'h1;
         mem[2321] = -3'h1;
         mem[2322] = -3'h1;
         mem[2323] = -3'h1;
         mem[2324] = -3'h1;
         mem[2325] = -3'h1;
         mem[2326] = -3'h1;
         mem[2327] = -3'h1;
         mem[2328] = -3'h1;
         mem[2329] = -3'h1;
         mem[2330] = -3'h1;
         mem[2331] = -3'h1;
         mem[2332] = -3'h1;
         mem[2333] = -3'h1;
         mem[2334] = -3'h1;
         mem[2335] = -3'h1;
         mem[2336] = -3'h1;
         mem[2337] = -3'h1;
         mem[2338] = -3'h1;
         mem[2339] = -3'h1;
         mem[2340] = -3'h1;
         mem[2341] = -3'h1;
         mem[2342] = -3'h1;
         mem[2343] = -3'h1;
         mem[2344] = -3'h1;
         mem[2345] = -3'h1;
         mem[2346] = -3'h1;
         mem[2347] = -3'h1;
         mem[2348] = -3'h1;
         mem[2349] = -3'h1;
         mem[2350] = -3'h1;
         mem[2351] = -3'h1;
         mem[2352] = -3'h1;
         mem[2353] = -3'h1;
         mem[2354] = -3'h1;
         mem[2355] = -3'h1;
         mem[2356] = -3'h1;
         mem[2357] = -3'h1;
         mem[2358] = -3'h1;
         mem[2359] = -3'h1;
         mem[2360] = -3'h1;
         mem[2361] = -3'h1;
         mem[2362] = -3'h1;
         mem[2363] = -3'h1;
         mem[2364] = -3'h1;
         mem[2365] = -3'h1;
         mem[2366] = -3'h1;
         mem[2367] = -3'h1;
         mem[2368] = -3'h1;
         mem[2369] = -3'h1;
         mem[2370] = -3'h1;
         mem[2371] = -3'h1;
         mem[2372] = -3'h1;
         mem[2373] = -3'h1;
         mem[2374] = -3'h1;
         mem[2375] = -3'h1;
         mem[2376] = -3'h1;
         mem[2377] = -3'h1;
         mem[2378] = -3'h1;
         mem[2379] = -3'h1;
         mem[2380] = -3'h1;
         mem[2381] = -3'h1;
         mem[2382] = -3'h1;
         mem[2383] = -3'h1;
         mem[2384] = -3'h1;
         mem[2385] = -3'h1;
         mem[2386] = -3'h1;
         mem[2387] = -3'h1;
         mem[2388] = -3'h1;
         mem[2389] = -3'h1;
         mem[2390] = -3'h1;
         mem[2391] = -3'h1;
         mem[2392] = -3'h1;
         mem[2393] = -3'h1;
         mem[2394] = -3'h1;
         mem[2395] = -3'h1;
         mem[2396] = -3'h1;
         mem[2397] = -3'h1;
         mem[2398] = -3'h1;
         mem[2399] = -3'h1;
         mem[2400] = -3'h1;
         mem[2401] = -3'h1;
         mem[2402] = -3'h1;
         mem[2403] = -3'h1;
         mem[2404] = -3'h1;
         mem[2405] = -3'h1;
         mem[2406] = -3'h1;
         mem[2407] = -3'h1;
         mem[2408] = -3'h1;
         mem[2409] = -3'h1;
         mem[2410] = -3'h1;
         mem[2411] = -3'h1;
         mem[2412] = -3'h1;
         mem[2413] = -3'h1;
         mem[2414] = -3'h1;
         mem[2415] = -3'h1;
         mem[2416] = -3'h1;
         mem[2417] = -3'h1;
         mem[2418] = -3'h1;
         mem[2419] = -3'h1;
         mem[2420] = -3'h1;
         mem[2421] = -3'h1;
         mem[2422] = -3'h1;
         mem[2423] = -3'h1;
         mem[2424] = -3'h1;
         mem[2425] = -3'h1;
         mem[2426] = -3'h1;
         mem[2427] = -3'h1;
         mem[2428] = -3'h1;
         mem[2429] = -3'h1;
         mem[2430] = -3'h1;
         mem[2431] = -3'h1;
         mem[2432] = -3'h1;
         mem[2433] = -3'h1;
         mem[2434] = -3'h1;
         mem[2435] = -3'h1;
         mem[2436] = -3'h1;
         mem[2437] = -3'h1;
         mem[2438] = -3'h1;
         mem[2439] = -3'h1;
         mem[2440] = -3'h1;
         mem[2441] = -3'h1;
         mem[2442] = -3'h1;
         mem[2443] = -3'h1;
         mem[2444] = -3'h1;
         mem[2445] = -3'h1;
         mem[2446] = -3'h1;
         mem[2447] = -3'h1;
         mem[2448] = -3'h1;
         mem[2449] = -3'h1;
         mem[2450] = -3'h1;
         mem[2451] = -3'h1;
         mem[2452] = -3'h1;
         mem[2453] = -3'h1;
         mem[2454] = -3'h1;
         mem[2455] = -3'h1;
         mem[2456] = -3'h1;
         mem[2457] = -3'h1;
         mem[2458] = -3'h1;
         mem[2459] = -3'h1;
         mem[2460] = -3'h1;
         mem[2461] = -3'h1;
         mem[2462] = -3'h1;
         mem[2463] = -3'h1;
         mem[2464] = -3'h1;
         mem[2465] = -3'h1;
         mem[2466] = -3'h1;
         mem[2467] = -3'h1;
         mem[2468] = -3'h1;
         mem[2469] = -3'h1;
         mem[2470] = -3'h1;
         mem[2471] = -3'h1;
         mem[2472] = -3'h1;
         mem[2473] = -3'h1;
         mem[2474] = -3'h1;
         mem[2475] = -3'h1;
         mem[2476] = -3'h1;
         mem[2477] = -3'h1;
         mem[2478] = -3'h1;
         mem[2479] = -3'h1;
         mem[2480] = -3'h1;
         mem[2481] = -3'h1;
         mem[2482] = -3'h1;
         mem[2483] = -3'h1;
         mem[2484] = -3'h1;
         mem[2485] = -3'h1;
         mem[2486] = -3'h1;
         mem[2487] = -3'h1;
         mem[2488] = -3'h1;
         mem[2489] = -3'h1;
         mem[2490] = -3'h1;
         mem[2491] = -3'h1;
         mem[2492] = -3'h1;
         mem[2493] = -3'h1;
         mem[2494] = -3'h1;
         mem[2495] = -3'h1;
         mem[2496] = -3'h1;
         mem[2497] = -3'h1;
         mem[2498] = -3'h1;
         mem[2499] = -3'h1;
         mem[2500] = -3'h1;
         mem[2501] = -3'h1;
         mem[2502] = -3'h1;
         mem[2503] = -3'h1;
         mem[2504] = -3'h1;
         mem[2505] = -3'h1;
         mem[2506] = -3'h1;
         mem[2507] = -3'h1;
         mem[2508] = -3'h1;
         mem[2509] = -3'h1;
         mem[2510] = -3'h1;
         mem[2511] = -3'h1;
         mem[2512] = -3'h1;
         mem[2513] = -3'h1;
         mem[2514] = -3'h1;
         mem[2515] = -3'h1;
         mem[2516] = -3'h1;
         mem[2517] = -3'h1;
         mem[2518] = -3'h1;
         mem[2519] = -3'h1;
         mem[2520] = -3'h1;
         mem[2521] = -3'h1;
         mem[2522] = -3'h1;
         mem[2523] = -3'h1;
         mem[2524] = -3'h1;
         mem[2525] = -3'h1;
         mem[2526] = -3'h1;
         mem[2527] = -3'h1;
         mem[2528] = -3'h1;
         mem[2529] = -3'h1;
         mem[2530] = -3'h1;
         mem[2531] = -3'h1;
         mem[2532] = -3'h1;
         mem[2533] = -3'h1;
         mem[2534] = -3'h1;
         mem[2535] = -3'h1;
         mem[2536] = -3'h1;
         mem[2537] = -3'h1;
         mem[2538] = -3'h1;
         mem[2539] = -3'h1;
         mem[2540] = -3'h1;
         mem[2541] = -3'h1;
         mem[2542] = -3'h1;
         mem[2543] = -3'h1;
         mem[2544] = -3'h1;
         mem[2545] = -3'h1;
         mem[2546] = -3'h1;
         mem[2547] = -3'h1;
         mem[2548] = -3'h1;
         mem[2549] = -3'h1;
         mem[2550] = -3'h1;
         mem[2551] = -3'h1;
         mem[2552] = -3'h1;
         mem[2553] = -3'h1;
         mem[2554] = -3'h1;
         mem[2555] = -3'h1;
         mem[2556] = -3'h1;
         mem[2557] = -3'h1;
         mem[2558] = -3'h1;
         mem[2559] = -3'h1;
         mem[2560] = -3'h1;
         mem[2561] = -3'h1;
         mem[2562] = -3'h1;
         mem[2563] = -3'h1;
         mem[2564] = -3'h1;
         mem[2565] = -3'h1;
         mem[2566] = -3'h1;
         mem[2567] = -3'h1;
         mem[2568] = -3'h1;
         mem[2569] = -3'h1;
         mem[2570] = -3'h1;
         mem[2571] = -3'h1;
         mem[2572] = -3'h1;
         mem[2573] = -3'h1;
         mem[2574] = -3'h1;
         mem[2575] = -3'h1;
         mem[2576] = -3'h1;
         mem[2577] = -3'h1;
         mem[2578] = -3'h1;
         mem[2579] = -3'h1;
         mem[2580] = -3'h1;
         mem[2581] = -3'h1;
         mem[2582] = -3'h1;
         mem[2583] = -3'h1;
         mem[2584] = -3'h1;
         mem[2585] = -3'h1;
         mem[2586] = -3'h1;
         mem[2587] = -3'h1;
         mem[2588] = -3'h1;
         mem[2589] = -3'h1;
         mem[2590] = -3'h1;
         mem[2591] = -3'h1;
         mem[2592] = -3'h1;
         mem[2593] = -3'h1;
         mem[2594] = -3'h1;
         mem[2595] = -3'h1;
         mem[2596] = -3'h1;
         mem[2597] = -3'h1;
         mem[2598] = -3'h1;
         mem[2599] = -3'h1;
         mem[2600] = -3'h1;
         mem[2601] = -3'h1;
         mem[2602] = -3'h1;
         mem[2603] = -3'h1;
         mem[2604] = -3'h1;
         mem[2605] = -3'h1;
         mem[2606] = -3'h1;
         mem[2607] = -3'h1;
         mem[2608] = -3'h1;
         mem[2609] = -3'h1;
         mem[2610] = -3'h1;
         mem[2611] = -3'h1;
         mem[2612] = -3'h1;
         mem[2613] = -3'h1;
         mem[2614] = -3'h1;
         mem[2615] = -3'h1;
         mem[2616] = -3'h1;
         mem[2617] = -3'h1;
         mem[2618] = -3'h1;
         mem[2619] = -3'h1;
         mem[2620] = -3'h1;
         mem[2621] = -3'h1;
         mem[2622] = -3'h1;
         mem[2623] = -3'h1;
         mem[2624] = -3'h1;
         mem[2625] = -3'h1;
         mem[2626] = -3'h1;
         mem[2627] = -3'h1;
         mem[2628] = -3'h1;
         mem[2629] = -3'h1;
         mem[2630] = -3'h1;
         mem[2631] = -3'h1;
         mem[2632] = -3'h1;
         mem[2633] = -3'h1;
         mem[2634] = -3'h1;
         mem[2635] = -3'h1;
         mem[2636] = -3'h1;
         mem[2637] = -3'h1;
         mem[2638] = -3'h1;
         mem[2639] = -3'h1;
         mem[2640] = -3'h1;
         mem[2641] = -3'h1;
         mem[2642] = -3'h1;
         mem[2643] = -3'h1;
         mem[2644] = -3'h1;
         mem[2645] = -3'h1;
         mem[2646] = -3'h1;
         mem[2647] = -3'h1;
         mem[2648] = -3'h1;
         mem[2649] = -3'h1;
         mem[2650] = -3'h1;
         mem[2651] = -3'h1;
         mem[2652] = -3'h1;
         mem[2653] = -3'h1;
         mem[2654] = -3'h1;
         mem[2655] = -3'h1;
         mem[2656] = -3'h1;
         mem[2657] = -3'h1;
         mem[2658] = -3'h1;
         mem[2659] = -3'h1;
         mem[2660] = -3'h1;
         mem[2661] = -3'h1;
         mem[2662] = -3'h1;
         mem[2663] = -3'h1;
         mem[2664] = -3'h1;
         mem[2665] = -3'h1;
         mem[2666] = -3'h1;
         mem[2667] = -3'h1;
         mem[2668] = -3'h1;
         mem[2669] = -3'h1;
         mem[2670] = -3'h1;
         mem[2671] = -3'h1;
         mem[2672] = -3'h1;
         mem[2673] = -3'h1;
         mem[2674] = -3'h1;
         mem[2675] = -3'h1;
         mem[2676] = -3'h1;
         mem[2677] = -3'h1;
         mem[2678] = -3'h1;
         mem[2679] = -3'h1;
         mem[2680] = -3'h1;
         mem[2681] = -3'h1;
         mem[2682] = -3'h1;
         mem[2683] = -3'h1;
         mem[2684] = -3'h1;
         mem[2685] = -3'h1;
         mem[2686] = -3'h1;
         mem[2687] = -3'h1;
         mem[2688] = -3'h1;
         mem[2689] = -3'h1;
         mem[2690] = -3'h1;
         mem[2691] = -3'h1;
         mem[2692] = -3'h1;
         mem[2693] = -3'h1;
         mem[2694] = -3'h1;
         mem[2695] = -3'h1;
         mem[2696] = -3'h1;
         mem[2697] = -3'h1;
         mem[2698] = -3'h1;
         mem[2699] = -3'h1;
         mem[2700] = -3'h1;
         mem[2701] = -3'h1;
         mem[2702] = -3'h1;
         mem[2703] = -3'h1;
         mem[2704] = -3'h1;
         mem[2705] = -3'h1;
         mem[2706] = -3'h1;
         mem[2707] = -3'h1;
         mem[2708] = -3'h1;
         mem[2709] = -3'h1;
         mem[2710] = -3'h1;
         mem[2711] = -3'h1;
         mem[2712] = -3'h1;
         mem[2713] = -3'h1;
         mem[2714] = -3'h1;
         mem[2715] = -3'h1;
         mem[2716] = -3'h1;
         mem[2717] = -3'h1;
         mem[2718] = -3'h1;
         mem[2719] = -3'h1;
         mem[2720] = -3'h1;
         mem[2721] = -3'h1;
         mem[2722] = -3'h1;
         mem[2723] = -3'h1;
         mem[2724] = -3'h1;
         mem[2725] = -3'h1;
         mem[2726] = -3'h1;
         mem[2727] = -3'h1;
         mem[2728] = -3'h1;
         mem[2729] = -3'h1;
         mem[2730] = -3'h1;
         mem[2731] = -3'h1;
         mem[2732] = -3'h1;
         mem[2733] = -3'h1;
         mem[2734] = -3'h1;
         mem[2735] = -3'h1;
         mem[2736] = -3'h1;
         mem[2737] = -3'h1;
         mem[2738] = -3'h1;
         mem[2739] = -3'h1;
         mem[2740] = -3'h1;
         mem[2741] = -3'h1;
         mem[2742] = -3'h1;
         mem[2743] = -3'h1;
         mem[2744] = -3'h1;
         mem[2745] = -3'h1;
         mem[2746] = -3'h1;
         mem[2747] = -3'h1;
         mem[2748] = -3'h1;
         mem[2749] = -3'h1;
         mem[2750] = -3'h1;
         mem[2751] = -3'h1;
         mem[2752] = -3'h1;
         mem[2753] = -3'h1;
         mem[2754] = -3'h1;
         mem[2755] = -3'h1;
         mem[2756] = -3'h1;
         mem[2757] = -3'h1;
         mem[2758] = -3'h1;
         mem[2759] = -3'h1;
         mem[2760] = -3'h1;
         mem[2761] = -3'h1;
         mem[2762] = -3'h1;
         mem[2763] = -3'h1;
         mem[2764] = -3'h1;
         mem[2765] = -3'h1;
         mem[2766] = -3'h1;
         mem[2767] = -3'h1;
         mem[2768] = -3'h1;
         mem[2769] = -3'h1;
         mem[2770] = -3'h1;
         mem[2771] = -3'h1;
         mem[2772] = -3'h1;
         mem[2773] = -3'h1;
         mem[2774] = -3'h1;
         mem[2775] = -3'h1;
         mem[2776] = -3'h1;
         mem[2777] = -3'h1;
         mem[2778] = -3'h1;
         mem[2779] = -3'h1;
         mem[2780] = -3'h1;
         mem[2781] = -3'h1;
         mem[2782] = -3'h1;
         mem[2783] = -3'h1;
         mem[2784] = -3'h1;
         mem[2785] = -3'h1;
         mem[2786] = -3'h1;
         mem[2787] = -3'h1;
         mem[2788] = -3'h1;
         mem[2789] = -3'h1;
         mem[2790] = -3'h1;
         mem[2791] = -3'h1;
         mem[2792] = -3'h1;
         mem[2793] = -3'h1;
         mem[2794] = -3'h1;
         mem[2795] = -3'h1;
         mem[2796] = -3'h1;
         mem[2797] = -3'h1;
         mem[2798] = -3'h1;
         mem[2799] = -3'h1;
         mem[2800] = -3'h1;
         mem[2801] = -3'h1;
         mem[2802] = -3'h1;
         mem[2803] = -3'h1;
         mem[2804] = -3'h1;
         mem[2805] = -3'h1;
         mem[2806] = -3'h1;
         mem[2807] = -3'h1;
         mem[2808] = -3'h1;
         mem[2809] = -3'h1;
         mem[2810] = -3'h1;
         mem[2811] = -3'h1;
         mem[2812] = -3'h1;
         mem[2813] = -3'h1;
         mem[2814] = -3'h1;
         mem[2815] = -3'h1;
         mem[2816] = -3'h1;
         mem[2817] = -3'h1;
         mem[2818] = -3'h1;
         mem[2819] = -3'h1;
         mem[2820] = -3'h1;
         mem[2821] = -3'h1;
         mem[2822] = -3'h1;
         mem[2823] = -3'h1;
         mem[2824] = -3'h1;
         mem[2825] = -3'h1;
         mem[2826] = -3'h1;
         mem[2827] = -3'h1;
         mem[2828] = -3'h1;
         mem[2829] = -3'h1;
         mem[2830] = -3'h1;
         mem[2831] = -3'h1;
         mem[2832] = -3'h1;
         mem[2833] = -3'h1;
         mem[2834] = -3'h1;
         mem[2835] = -3'h1;
         mem[2836] = -3'h1;
         mem[2837] = -3'h1;
         mem[2838] = -3'h1;
         mem[2839] = -3'h1;
         mem[2840] = -3'h1;
         mem[2841] = -3'h1;
         mem[2842] = -3'h1;
         mem[2843] = -3'h1;
         mem[2844] = -3'h1;
         mem[2845] = -3'h1;
         mem[2846] = -3'h1;
         mem[2847] = -3'h1;
         mem[2848] = -3'h1;
         mem[2849] = -3'h1;
         mem[2850] = -3'h1;
         mem[2851] = -3'h1;
         mem[2852] = -3'h1;
         mem[2853] = -3'h1;
         mem[2854] = -3'h1;
         mem[2855] = -3'h1;
         mem[2856] = -3'h1;
         mem[2857] = -3'h1;
         mem[2858] = -3'h1;
         mem[2859] = -3'h1;
         mem[2860] = -3'h1;
         mem[2861] = -3'h1;
         mem[2862] = -3'h1;
         mem[2863] = -3'h1;
         mem[2864] = -3'h1;
         mem[2865] = -3'h1;
         mem[2866] = -3'h1;
         mem[2867] = -3'h1;
         mem[2868] = -3'h1;
         mem[2869] = -3'h1;
         mem[2870] = -3'h1;
         mem[2871] = -3'h1;
         mem[2872] = -3'h1;
         mem[2873] = -3'h1;
         mem[2874] = -3'h1;
         mem[2875] = -3'h1;
         mem[2876] = -3'h1;
         mem[2877] = -3'h1;
         mem[2878] = -3'h1;
         mem[2879] = -3'h1;
         mem[2880] = -3'h1;
         mem[2881] = -3'h1;
         mem[2882] = -3'h1;
         mem[2883] = -3'h1;
         mem[2884] = -3'h1;
         mem[2885] = -3'h1;
         mem[2886] = -3'h1;
         mem[2887] = -3'h1;
         mem[2888] = -3'h1;
         mem[2889] = -3'h1;
         mem[2890] = -3'h1;
         mem[2891] = -3'h1;
         mem[2892] = -3'h1;
         mem[2893] = -3'h1;
         mem[2894] = -3'h1;
         mem[2895] = -3'h1;
         mem[2896] = -3'h1;
         mem[2897] = -3'h1;
         mem[2898] = -3'h1;
         mem[2899] = -3'h1;
         mem[2900] = -3'h1;
         mem[2901] = -3'h1;
         mem[2902] = -3'h1;
         mem[2903] = -3'h1;
         mem[2904] = -3'h1;
         mem[2905] = -3'h1;
         mem[2906] = -3'h1;
         mem[2907] = -3'h1;
         mem[2908] = -3'h1;
         mem[2909] = -3'h1;
         mem[2910] = -3'h1;
         mem[2911] = -3'h1;
         mem[2912] = -3'h1;
     end

endmodule: weights0_rom
