module featureThreshold_rom
  #(
     W_DATA = 13,
     DEPTH = 2913,
     W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input ena,
     input [W_ADDR-1:0] addra,
     output [W_DATA-1:0] doa
    );

     (* rom_style = "block" *)


     logic [W_DATA-1:0] mem [DEPTH-1:0];

     always_ff @(posedge clk)
        begin
           if(ena)
              doa = mem[addra];
        end

     initial begin
         mem[0] = -13'h0081;
         mem[1] =  13'h0032;
         mem[2] =  13'h0059;
         mem[3] =  13'h0017;
         mem[4] =  13'h003d;
         mem[5] =  13'h0197;
         mem[6] =  13'h000b;
         mem[7] = -13'h004d;
         mem[8] =  13'h0018;
         mem[9] = -13'h0056;
         mem[10] =  13'h0053;
         mem[11] =  13'h0057;
         mem[12] =  13'h0177;
         mem[13] =  13'h0094;
         mem[14] = -13'h004e;
         mem[15] =  13'h0021;
         mem[16] =  13'h004b;
         mem[17] = -13'h001c;
         mem[18] = -13'h0028;
         mem[19] =  13'h0040;
         mem[20] = -13'h0054;
         mem[21] = -13'h0233;
         mem[22] =  13'h003a;
         mem[23] =  13'h0029;
         mem[24] =  13'h0176;
         mem[25] =  13'h011d;
         mem[26] =  13'h0081;
         mem[27] =  13'h003a;
         mem[28] =  13'h003b;
         mem[29] = -13'h000c;
         mem[30] =  13'h0086;
         mem[31] = -13'h001d;
         mem[32] =  13'h00ce;
         mem[33] =  13'h00c0;
         mem[34] = -13'h011c;
         mem[35] = -13'h00c8;
         mem[36] =  13'h015b;
         mem[37] = -13'h0007;
         mem[38] =  13'h01d9;
         mem[39] = -13'h00d2;
         mem[40] = -13'h00ae;
         mem[41] =  13'h05f2;
         mem[42] =  13'h004f;
         mem[43] =  13'h0047;
         mem[44] =  13'h00a2;
         mem[45] = -13'h0025;
         mem[46] =  13'h0007;
         mem[47] =  13'h007b;
         mem[48] = -13'h0142;
         mem[49] =  13'h0008;
         mem[50] =  13'h006e;
         mem[51] = -13'h00b8;
         mem[52] = -13'h010d;
         mem[53] =  13'h0040;
         mem[54] =  13'h0254;
         mem[55] =  13'h0019;
         mem[56] =  13'h001b;
         mem[57] =  13'h004b;
         mem[58] =  13'h0051;
         mem[59] = -13'h0470;
         mem[60] =  13'h0025;
         mem[61] = -13'h009a;
         mem[62] =  13'h004b;
         mem[63] = -13'h002d;
         mem[64] =  13'h008a;
         mem[65] = -13'h0092;
         mem[66] = -13'h002e;
         mem[67] = -13'h010b;
         mem[68] = -13'h00ad;
         mem[69] =  13'h0007;
         mem[70] = -13'h0211;
         mem[71] =  13'h005d;
         mem[72] = -13'h008b;
         mem[73] =  13'h006b;
         mem[74] =  13'h005b;
         mem[75] = -13'h0017;
         mem[76] =  13'h00b2;
         mem[77] =  13'h00ea;
         mem[78] =  13'h0009;
         mem[79] =  13'h0035;
         mem[80] = -13'h006c;
         mem[81] = -13'h0017;
         mem[82] = -13'h0043;
         mem[83] = -13'h0117;
         mem[84] =  13'h00a3;
         mem[85] =  13'h0302;
         mem[86] =  13'h013f;
         mem[87] =  13'h0000;
         mem[88] =  13'h015c;
         mem[89] =  13'h0024;
         mem[90] =  13'h0024;
         mem[91] = -13'h0060;
         mem[92] =  13'h001c;
         mem[93] =  13'h008a;
         mem[94] = -13'h000d;
         mem[95] =  13'h0077;
         mem[96] = -13'h0022;
         mem[97] = -13'h002c;
         mem[98] = -13'h0064;
         mem[99] =  13'h000f;
         mem[100] = -13'h0032;
         mem[101] = -13'h0013;
         mem[102] =  13'h013a;
         mem[103] =  13'h0075;
         mem[104] =  13'h0050;
         mem[105] = -13'h0077;
         mem[106] = -13'h0077;
         mem[107] =  13'h0050;
         mem[108] =  13'h0011;
         mem[109] = -13'h0091;
         mem[110] = -13'h0042;
         mem[111] = -13'h005a;
         mem[112] = -13'h005d;
         mem[113] =  13'h0044;
         mem[114] = -13'h0036;
         mem[115] = -13'h008a;
         mem[116] =  13'h0045;
         mem[117] =  13'h000d;
         mem[118] =  13'h0156;
         mem[119] =  13'h0420;
         mem[120] = -13'h0095;
         mem[121] = -13'h0043;
         mem[122] = -13'h000f;
         mem[123] = -13'h001a;
         mem[124] = -13'h000f;
         mem[125] = -13'h00ba;
         mem[126] = -13'h0062;
         mem[127] = -13'h013d;
         mem[128] =  13'h0060;
         mem[129] = -13'h000a;
         mem[130] =  13'h01eb;
         mem[131] =  13'h0009;
         mem[132] =  13'h011d;
         mem[133] = -13'h00bf;
         mem[134] = -13'h00cd;
         mem[135] =  13'h007b;
         mem[136] =  13'h0175;
         mem[137] =  13'h0034;
         mem[138] =  13'h0041;
         mem[139] =  13'h0009;
         mem[140] =  13'h0082;
         mem[141] =  13'h000b;
         mem[142] = -13'h0031;
         mem[143] =  13'h0057;
         mem[144] =  13'h007c;
         mem[145] = -13'h00b8;
         mem[146] = -13'h0125;
         mem[147] =  13'h00f2;
         mem[148] =  13'h001b;
         mem[149] =  13'h00a8;
         mem[150] = -13'h0003;
         mem[151] = -13'h007c;
         mem[152] = -13'h0034;
         mem[153] =  13'h0099;
         mem[154] =  13'h0064;
         mem[155] =  13'h00e9;
         mem[156] = -13'h0042;
         mem[157] = -13'h02d2;
         mem[158] =  13'h02d1;
         mem[159] = -13'h001e;
         mem[160] =  13'h00f9;
         mem[161] = -13'h0077;
         mem[162] = -13'h00ba;
         mem[163] =  13'h0098;
         mem[164] = -13'h0063;
         mem[165] = -13'h00f4;
         mem[166] = -13'h007b;
         mem[167] =  13'h001e;
         mem[168] = -13'h0008;
         mem[169] =  13'h0055;
         mem[170] = -13'h001b;
         mem[171] =  13'h004c;
         mem[172] = -13'h00b5;
         mem[173] =  13'h005d;
         mem[174] = -13'h0004;
         mem[175] =  13'h0046;
         mem[176] = -13'h008d;
         mem[177] =  13'h0112;
         mem[178] =  13'h03cd;
         mem[179] = -13'h0034;
         mem[180] =  13'h002b;
         mem[181] =  13'h0045;
         mem[182] = -13'h001d;
         mem[183] =  13'h002b;
         mem[184] =  13'h0019;
         mem[185] =  13'h0035;
         mem[186] =  13'h000c;
         mem[187] = -13'h01bf;
         mem[188] =  13'h0021;
         mem[189] =  13'h0080;
         mem[190] =  13'h0082;
         mem[191] =  13'h001b;
         mem[192] =  13'h006b;
         mem[193] =  13'h0034;
         mem[194] =  13'h006b;
         mem[195] = -13'h003d;
         mem[196] = -13'h009f;
         mem[197] = -13'h0017;
         mem[198] = -13'h0006;
         mem[199] = -13'h0074;
         mem[200] =  13'h010f;
         mem[201] =  13'h0024;
         mem[202] =  13'h002e;
         mem[203] = -13'h000b;
         mem[204] =  13'h002e;
         mem[205] =  13'h001d;
         mem[206] =  13'h0082;
         mem[207] =  13'h0067;
         mem[208] =  13'h001e;
         mem[209] =  13'h0086;
         mem[210] = -13'h000b;
         mem[211] = -13'h009b;
         mem[212] = -13'h009f;
         mem[213] =  13'h000b;
         mem[214] = -13'h00dd;
         mem[215] = -13'h0022;
         mem[216] =  13'h008a;
         mem[217] = -13'h01cc;
         mem[218] = -13'h002a;
         mem[219] = -13'h0014;
         mem[220] = -13'h0026;
         mem[221] = -13'h0030;
         mem[222] = -13'h005f;
         mem[223] =  13'h0045;
         mem[224] = -13'h0062;
         mem[225] = -13'h0097;
         mem[226] = -13'h00fc;
         mem[227] =  13'h0058;
         mem[228] = -13'h000f;
         mem[229] =  13'h00b7;
         mem[230] =  13'h00ea;
         mem[231] = -13'h002e;
         mem[232] = -13'h0031;
         mem[233] =  13'h005c;
         mem[234] = -13'h0051;
         mem[235] =  13'h0041;
         mem[236] = -13'h0025;
         mem[237] = -13'h0012;
         mem[238] =  13'h0209;
         mem[239] =  13'h00c3;
         mem[240] =  13'h00db;
         mem[241] = -13'h00a2;
         mem[242] = -13'h0113;
         mem[243] =  13'h0222;
         mem[244] = -13'h0358;
         mem[245] = -13'h010c;
         mem[246] =  13'h00fd;
         mem[247] = -13'h0068;
         mem[248] = -13'h008e;
         mem[249] = -13'h004a;
         mem[250] =  13'h003d;
         mem[251] =  13'h00bd;
         mem[252] =  13'h003f;
         mem[253] =  13'h0034;
         mem[254] =  13'h00c9;
         mem[255] =  13'h0033;
         mem[256] = -13'h004c;
         mem[257] =  13'h00ab;
         mem[258] = -13'h00d2;
         mem[259] = -13'h0122;
         mem[260] =  13'h0044;
         mem[261] = -13'h0019;
         mem[262] = -13'h00a1;
         mem[263] =  13'h0000;
         mem[264] = -13'h005b;
         mem[265] =  13'h0007;
         mem[266] =  13'h0004;
         mem[267] =  13'h00a0;
         mem[268] =  13'h00fe;
         mem[269] =  13'h0008;
         mem[270] =  13'h0003;
         mem[271] = -13'h001c;
         mem[272] = -13'h0061;
         mem[273] = -13'h01a4;
         mem[274] = -13'h0027;
         mem[275] =  13'h00a3;
         mem[276] = -13'h0035;
         mem[277] = -13'h00cf;
         mem[278] =  13'h0066;
         mem[279] = -13'h001f;
         mem[280] =  13'h00af;
         mem[281] =  13'h0000;
         mem[282] =  13'h0025;
         mem[283] =  13'h002d;
         mem[284] = -13'h00d6;
         mem[285] = -13'h03ae;
         mem[286] = -13'h0043;
         mem[287] = -13'h0046;
         mem[288] = -13'h0096;
         mem[289] = -13'h002a;
         mem[290] = -13'h0038;
         mem[291] =  13'h0078;
         mem[292] =  13'h0062;
         mem[293] =  13'h0019;
         mem[294] = -13'h005b;
         mem[295] = -13'h001c;
         mem[296] = -13'h00a6;
         mem[297] = -13'h0064;
         mem[298] =  13'h000a;
         mem[299] = -13'h0050;
         mem[300] = -13'h0079;
         mem[301] = -13'h003d;
         mem[302] = -13'h00f8;
         mem[303] = -13'h0034;
         mem[304] = -13'h0052;
         mem[305] = -13'h007d;
         mem[306] = -13'h0054;
         mem[307] = -13'h0007;
         mem[308] = -13'h0080;
         mem[309] =  13'h004d;
         mem[310] =  13'h0019;
         mem[311] = -13'h0029;
         mem[312] = -13'h0005;
         mem[313] = -13'h0010;
         mem[314] = -13'h00b4;
         mem[315] = -13'h00f8;
         mem[316] = -13'h0086;
         mem[317] = -13'h025b;
         mem[318] = -13'h0030;
         mem[319] =  13'h0252;
         mem[320] =  13'h00d2;
         mem[321] =  13'h000c;
         mem[322] = -13'h00b2;
         mem[323] =  13'h0210;
         mem[324] = -13'h0175;
         mem[325] =  13'h003a;
         mem[326] =  13'h0086;
         mem[327] =  13'h0033;
         mem[328] =  13'h003c;
         mem[329] = -13'h0089;
         mem[330] =  13'h0247;
         mem[331] = -13'h0019;
         mem[332] =  13'h004a;
         mem[333] =  13'h0066;
         mem[334] =  13'h00be;
         mem[335] = -13'h0024;
         mem[336] =  13'h00a7;
         mem[337] = -13'h008c;
         mem[338] = -13'h00a2;
         mem[339] =  13'h000a;
         mem[340] =  13'h0070;
         mem[341] =  13'h008f;
         mem[342] =  13'h0012;
         mem[343] =  13'h000b;
         mem[344] =  13'h0090;
         mem[345] =  13'h006a;
         mem[346] = -13'h0040;
         mem[347] = -13'h001f;
         mem[348] =  13'h0055;
         mem[349] =  13'h00f5;
         mem[350] =  13'h009f;
         mem[351] =  13'h0058;
         mem[352] = -13'h0070;
         mem[353] =  13'h002a;
         mem[354] =  13'h0065;
         mem[355] = -13'h0041;
         mem[356] =  13'h00c7;
         mem[357] =  13'h0005;
         mem[358] = -13'h0168;
         mem[359] =  13'h004b;
         mem[360] =  13'h0090;
         mem[361] = -13'h0343;
         mem[362] = -13'h0044;
         mem[363] =  13'h009a;
         mem[364] =  13'h0009;
         mem[365] = -13'h003c;
         mem[366] = -13'h00c5;
         mem[367] = -13'h0078;
         mem[368] = -13'h00bd;
         mem[369] = -13'h0072;
         mem[370] = -13'h0017;
         mem[371] = -13'h0029;
         mem[372] =  13'h002e;
         mem[373] =  13'h00d4;
         mem[374] =  13'h0088;
         mem[375] = -13'h003b;
         mem[376] = -13'h008c;
         mem[377] = -13'h014a;
         mem[378] = -13'h0003;
         mem[379] =  13'h018d;
         mem[380] =  13'h0095;
         mem[381] =  13'h00d3;
         mem[382] = -13'h0064;
         mem[383] =  13'h053c;
         mem[384] =  13'h001f;
         mem[385] =  13'h0296;
         mem[386] = -13'h0013;
         mem[387] = -13'h004b;
         mem[388] =  13'h013e;
         mem[389] =  13'h004d;
         mem[390] = -13'h0145;
         mem[391] = -13'h0116;
         mem[392] = -13'h0018;
         mem[393] =  13'h0082;
         mem[394] = -13'h007a;
         mem[395] = -13'h0149;
         mem[396] =  13'h000f;
         mem[397] =  13'h0089;
         mem[398] =  13'h0021;
         mem[399] =  13'h019d;
         mem[400] = -13'h0028;
         mem[401] =  13'h001d;
         mem[402] =  13'h0066;
         mem[403] =  13'h0477;
         mem[404] = -13'h00b5;
         mem[405] = -13'h0039;
         mem[406] =  13'h0234;
         mem[407] =  13'h008d;
         mem[408] =  13'h004c;
         mem[409] =  13'h0066;
         mem[410] =  13'h00ea;
         mem[411] =  13'h003d;
         mem[412] =  13'h0024;
         mem[413] =  13'h007c;
         mem[414] = -13'h00b4;
         mem[415] =  13'h004b;
         mem[416] =  13'h002b;
         mem[417] = -13'h00bc;
         mem[418] =  13'h0153;
         mem[419] = -13'h0024;
         mem[420] =  13'h00af;
         mem[421] = -13'h0023;
         mem[422] = -13'h0011;
         mem[423] =  13'h0021;
         mem[424] =  13'h018c;
         mem[425] = -13'h007d;
         mem[426] = -13'h00f9;
         mem[427] = -13'h009c;
         mem[428] = -13'h0027;
         mem[429] =  13'h00c8;
         mem[430] = -13'h00aa;
         mem[431] = -13'h0052;
         mem[432] = -13'h0004;
         mem[433] = -13'h0089;
         mem[434] =  13'h004f;
         mem[435] = -13'h0001;
         mem[436] = -13'h0001;
         mem[437] = -13'h017e;
         mem[438] = -13'h013e;
         mem[439] =  13'h0045;
         mem[440] = -13'h0057;
         mem[441] = -13'h0034;
         mem[442] =  13'h0020;
         mem[443] =  13'h01a5;
         mem[444] = -13'h0099;
         mem[445] =  13'h0068;
         mem[446] =  13'h0002;
         mem[447] = -13'h049e;
         mem[448] =  13'h0175;
         mem[449] =  13'h01ed;
         mem[450] = -13'h012e;
         mem[451] = -13'h0087;
         mem[452] = -13'h00b3;
         mem[453] =  13'h02e5;
         mem[454] = -13'h0030;
         mem[455] =  13'h0012;
         mem[456] =  13'h001c;
         mem[457] = -13'h0061;
         mem[458] = -13'h0113;
         mem[459] = -13'h010b;
         mem[460] =  13'h005d;
         mem[461] = -13'h004d;
         mem[462] = -13'h001c;
         mem[463] = -13'h00a4;
         mem[464] = -13'h00a6;
         mem[465] = -13'h0032;
         mem[466] = -13'h006f;
         mem[467] = -13'h0169;
         mem[468] = -13'h0020;
         mem[469] = -13'h00ab;
         mem[470] =  13'h00bb;
         mem[471] = -13'h0241;
         mem[472] = -13'h00f2;
         mem[473] =  13'h0011;
         mem[474] = -13'h0008;
         mem[475] =  13'h0467;
         mem[476] = -13'h006c;
         mem[477] =  13'h00a7;
         mem[478] =  13'h0016;
         mem[479] =  13'h0082;
         mem[480] = -13'h00a9;
         mem[481] = -13'h0189;
         mem[482] = -13'h002f;
         mem[483] =  13'h004b;
         mem[484] = -13'h008b;
         mem[485] = -13'h0064;
         mem[486] =  13'h00c8;
         mem[487] = -13'h0054;
         mem[488] = -13'h005e;
         mem[489] =  13'h0108;
         mem[490] =  13'h0033;
         mem[491] = -13'h0031;
         mem[492] = -13'h006c;
         mem[493] = -13'h0068;
         mem[494] =  13'h00a0;
         mem[495] = -13'h0018;
         mem[496] = -13'h008b;
         mem[497] =  13'h00a6;
         mem[498] =  13'h0068;
         mem[499] =  13'h0331;
         mem[500] =  13'h0032;
         mem[501] =  13'h00a0;
         mem[502] = -13'h007e;
         mem[503] = -13'h0091;
         mem[504] = -13'h00fc;
         mem[505] = -13'h0030;
         mem[506] =  13'h0112;
         mem[507] = -13'h0054;
         mem[508] = -13'h005b;
         mem[509] =  13'h0004;
         mem[510] =  13'h0092;
         mem[511] =  13'h007d;
         mem[512] =  13'h0016;
         mem[513] = -13'h0019;
         mem[514] = -13'h007c;
         mem[515] = -13'h0027;
         mem[516] = -13'h00e9;
         mem[517] =  13'h0010;
         mem[518] =  13'h008a;
         mem[519] = -13'h008d;
         mem[520] =  13'h00c0;
         mem[521] = -13'h0023;
         mem[522] =  13'h010c;
         mem[523] = -13'h00b4;
         mem[524] =  13'h0046;
         mem[525] =  13'h0087;
         mem[526] = -13'h0056;
         mem[527] =  13'h0079;
         mem[528] =  13'h00e2;
         mem[529] = -13'h0089;
         mem[530] =  13'h0050;
         mem[531] = -13'h0055;
         mem[532] =  13'h0085;
         mem[533] = -13'h002c;
         mem[534] = -13'h0028;
         mem[535] = -13'h000f;
         mem[536] = -13'h00ab;
         mem[537] = -13'h008c;
         mem[538] =  13'h0029;
         mem[539] = -13'h0170;
         mem[540] =  13'h006a;
         mem[541] = -13'h000f;
         mem[542] =  13'h0082;
         mem[543] =  13'h004f;
         mem[544] =  13'h0007;
         mem[545] = -13'h00b4;
         mem[546] = -13'h00b7;
         mem[547] = -13'h01b8;
         mem[548] = -13'h020e;
         mem[549] = -13'h00b7;
         mem[550] = -13'h00b4;
         mem[551] = -13'h01f6;
         mem[552] = -13'h0051;
         mem[553] = -13'h003f;
         mem[554] = -13'h00c8;
         mem[555] =  13'h00e5;
         mem[556] = -13'h0028;
         mem[557] =  13'h0037;
         mem[558] =  13'h001a;
         mem[559] =  13'h001d;
         mem[560] =  13'h0013;
         mem[561] =  13'h0027;
         mem[562] = -13'h0070;
         mem[563] = -13'h00a1;
         mem[564] = -13'h007d;
         mem[565] = -13'h0006;
         mem[566] =  13'h030d;
         mem[567] =  13'h0015;
         mem[568] =  13'h0062;
         mem[569] = -13'h006c;
         mem[570] =  13'h0016;
         mem[571] =  13'h00de;
         mem[572] =  13'h0000;
         mem[573] =  13'h003e;
         mem[574] =  13'h0045;
         mem[575] =  13'h007c;
         mem[576] =  13'h001a;
         mem[577] =  13'h0244;
         mem[578] =  13'h004f;
         mem[579] = -13'h0046;
         mem[580] = -13'h0019;
         mem[581] = -13'h0041;
         mem[582] = -13'h019e;
         mem[583] = -13'h001e;
         mem[584] =  13'h00b5;
         mem[585] = -13'h01dc;
         mem[586] =  13'h0013;
         mem[587] =  13'h005b;
         mem[588] = -13'h0031;
         mem[589] =  13'h00e5;
         mem[590] = -13'h0023;
         mem[591] =  13'h001b;
         mem[592] = -13'h004a;
         mem[593] = -13'h005d;
         mem[594] =  13'h0034;
         mem[595] = -13'h0038;
         mem[596] =  13'h0080;
         mem[597] =  13'h017d;
         mem[598] =  13'h006a;
         mem[599] =  13'h0043;
         mem[600] = -13'h0007;
         mem[601] = -13'h0024;
         mem[602] =  13'h005c;
         mem[603] = -13'h009a;
         mem[604] = -13'h0016;
         mem[605] = -13'h0061;
         mem[606] = -13'h006c;
         mem[607] =  13'h0032;
         mem[608] =  13'h018b;
         mem[609] = -13'h0070;
         mem[610] = -13'h0040;
         mem[611] = -13'h0008;
         mem[612] =  13'h0031;
         mem[613] = -13'h003f;
         mem[614] = -13'h0011;
         mem[615] = -13'h0056;
         mem[616] = -13'h0045;
         mem[617] = -13'h00a7;
         mem[618] = -13'h0021;
         mem[619] = -13'h004e;
         mem[620] = -13'h00b5;
         mem[621] = -13'h00ff;
         mem[622] = -13'h0004;
         mem[623] =  13'h0061;
         mem[624] =  13'h0057;
         mem[625] =  13'h0052;
         mem[626] = -13'h0075;
         mem[627] =  13'h000e;
         mem[628] =  13'h00e9;
         mem[629] = -13'h0180;
         mem[630] =  13'h0048;
         mem[631] =  13'h03a7;
         mem[632] = -13'h02ed;
         mem[633] = -13'h011e;
         mem[634] =  13'h003e;
         mem[635] =  13'h001b;
         mem[636] = -13'h0041;
         mem[637] =  13'h0035;
         mem[638] =  13'h0035;
         mem[639] = -13'h00a3;
         mem[640] =  13'h003d;
         mem[641] = -13'h0054;
         mem[642] = -13'h005b;
         mem[643] = -13'h0020;
         mem[644] =  13'h003e;
         mem[645] = -13'h0081;
         mem[646] = -13'h007e;
         mem[647] = -13'h003f;
         mem[648] =  13'h0090;
         mem[649] = -13'h0049;
         mem[650] = -13'h000d;
         mem[651] =  13'h0040;
         mem[652] =  13'h007a;
         mem[653] =  13'h000c;
         mem[654] =  13'h015b;
         mem[655] = -13'h00f0;
         mem[656] =  13'h00b7;
         mem[657] =  13'h00a5;
         mem[658] =  13'h009a;
         mem[659] =  13'h00f8;
         mem[660] = -13'h0051;
         mem[661] = -13'h02a7;
         mem[662] =  13'h011a;
         mem[663] =  13'h002e;
         mem[664] =  13'h0006;
         mem[665] =  13'h0146;
         mem[666] = -13'h00ea;
         mem[667] =  13'h001e;
         mem[668] = -13'h0049;
         mem[669] =  13'h0183;
         mem[670] =  13'h0016;
         mem[671] =  13'h001c;
         mem[672] =  13'h008d;
         mem[673] = -13'h00d4;
         mem[674] = -13'h011b;
         mem[675] = -13'h0016;
         mem[676] =  13'h0118;
         mem[677] = -13'h0112;
         mem[678] = -13'h0056;
         mem[679] =  13'h0053;
         mem[680] = -13'h00c0;
         mem[681] =  13'h0300;
         mem[682] = -13'h00b1;
         mem[683] =  13'h0051;
         mem[684] =  13'h0021;
         mem[685] =  13'h006f;
         mem[686] = -13'h0177;
         mem[687] = -13'h0033;
         mem[688] =  13'h003c;
         mem[689] =  13'h0077;
         mem[690] =  13'h0023;
         mem[691] = -13'h00e0;
         mem[692] = -13'h003c;
         mem[693] =  13'h0066;
         mem[694] =  13'h00be;
         mem[695] =  13'h0048;
         mem[696] =  13'h029c;
         mem[697] =  13'h0035;
         mem[698] = -13'h0040;
         mem[699] =  13'h0149;
         mem[700] =  13'h0090;
         mem[701] =  13'h0087;
         mem[702] =  13'h0031;
         mem[703] =  13'h00b0;
         mem[704] =  13'h007c;
         mem[705] =  13'h0091;
         mem[706] = -13'h003b;
         mem[707] =  13'h0033;
         mem[708] =  13'h0029;
         mem[709] =  13'h0076;
         mem[710] =  13'h0002;
         mem[711] =  13'h00c6;
         mem[712] =  13'h0084;
         mem[713] =  13'h0088;
         mem[714] =  13'h001a;
         mem[715] = -13'h0017;
         mem[716] =  13'h0034;
         mem[717] =  13'h0018;
         mem[718] =  13'h000a;
         mem[719] = -13'h0045;
         mem[720] =  13'h0073;
         mem[721] =  13'h002a;
         mem[722] =  13'h0028;
         mem[723] =  13'h006a;
         mem[724] = -13'h0068;
         mem[725] = -13'h000e;
         mem[726] =  13'h0025;
         mem[727] =  13'h0056;
         mem[728] = -13'h00d1;
         mem[729] = -13'h00ff;
         mem[730] = -13'h0087;
         mem[731] = -13'h0099;
         mem[732] =  13'h01fc;
         mem[733] = -13'h0024;
         mem[734] = -13'h00f5;
         mem[735] =  13'h0019;
         mem[736] = -13'h0048;
         mem[737] =  13'h0048;
         mem[738] =  13'h0015;
         mem[739] = -13'h002b;
         mem[740] =  13'h0357;
         mem[741] = -13'h006c;
         mem[742] =  13'h00f1;
         mem[743] = -13'h002f;
         mem[744] =  13'h00bc;
         mem[745] = -13'h005d;
         mem[746] = -13'h0021;
         mem[747] =  13'h000e;
         mem[748] =  13'h00ca;
         mem[749] =  13'h000e;
         mem[750] = -13'h007e;
         mem[751] =  13'h0162;
         mem[752] = -13'h022f;
         mem[753] = -13'h0017;
         mem[754] = -13'h0049;
         mem[755] = -13'h0051;
         mem[756] = -13'h00eb;
         mem[757] = -13'h0154;
         mem[758] = -13'h00dc;
         mem[759] = -13'h0022;
         mem[760] =  13'h00e2;
         mem[761] = -13'h0113;
         mem[762] = -13'h0061;
         mem[763] =  13'h0016;
         mem[764] =  13'h0057;
         mem[765] = -13'h0064;
         mem[766] = -13'h0050;
         mem[767] = -13'h00da;
         mem[768] =  13'h001d;
         mem[769] = -13'h005c;
         mem[770] = -13'h0151;
         mem[771] =  13'h0218;
         mem[772] =  13'h003a;
         mem[773] =  13'h001a;
         mem[774] = -13'h00bc;
         mem[775] =  13'h00ec;
         mem[776] = -13'h0018;
         mem[777] = -13'h00d5;
         mem[778] =  13'h00be;
         mem[779] =  13'h001e;
         mem[780] =  13'h0058;
         mem[781] = -13'h0049;
         mem[782] = -13'h0098;
         mem[783] = -13'h0001;
         mem[784] =  13'h0066;
         mem[785] =  13'h0026;
         mem[786] =  13'h0084;
         mem[787] = -13'h0019;
         mem[788] =  13'h00d2;
         mem[789] = -13'h006c;
         mem[790] = -13'h003f;
         mem[791] =  13'h004f;
         mem[792] =  13'h0089;
         mem[793] =  13'h0076;
         mem[794] =  13'h0000;
         mem[795] = -13'h00c9;
         mem[796] =  13'h0139;
         mem[797] =  13'h0061;
         mem[798] =  13'h000f;
         mem[799] = -13'h016e;
         mem[800] = -13'h003d;
         mem[801] = -13'h002d;
         mem[802] =  13'h0183;
         mem[803] =  13'h08ce;
         mem[804] =  13'h00a9;
         mem[805] =  13'h0065;
         mem[806] =  13'h00d0;
         mem[807] = -13'h0045;
         mem[808] = -13'h01f2;
         mem[809] = -13'h000e;
         mem[810] =  13'h01da;
         mem[811] =  13'h0097;
         mem[812] =  13'h002f;
         mem[813] = -13'h0052;
         mem[814] = -13'h0075;
         mem[815] = -13'h0017;
         mem[816] = -13'h00e3;
         mem[817] = -13'h003c;
         mem[818] = -13'h001d;
         mem[819] = -13'h00b8;
         mem[820] =  13'h0107;
         mem[821] = -13'h003c;
         mem[822] =  13'h00b8;
         mem[823] = -13'h0004;
         mem[824] =  13'h00ca;
         mem[825] =  13'h0077;
         mem[826] =  13'h008e;
         mem[827] = -13'h0019;
         mem[828] =  13'h003f;
         mem[829] =  13'h000b;
         mem[830] = -13'h00db;
         mem[831] = -13'h004e;
         mem[832] = -13'h00e2;
         mem[833] =  13'h00e6;
         mem[834] = -13'h0061;
         mem[835] =  13'h0007;
         mem[836] = -13'h009a;
         mem[837] = -13'h0062;
         mem[838] =  13'h0070;
         mem[839] =  13'h01d9;
         mem[840] = -13'h005b;
         mem[841] =  13'h0036;
         mem[842] = -13'h000f;
         mem[843] = -13'h000a;
         mem[844] =  13'h000d;
         mem[845] =  13'h009a;
         mem[846] = -13'h0038;
         mem[847] = -13'h000b;
         mem[848] = -13'h009d;
         mem[849] = -13'h008e;
         mem[850] =  13'h005f;
         mem[851] =  13'h008f;
         mem[852] = -13'h0036;
         mem[853] =  13'h0034;
         mem[854] =  13'h000e;
         mem[855] =  13'h019c;
         mem[856] =  13'h0000;
         mem[857] =  13'h002f;
         mem[858] = -13'h0093;
         mem[859] = -13'h0056;
         mem[860] =  13'h003c;
         mem[861] = -13'h0015;
         mem[862] =  13'h0060;
         mem[863] = -13'h0066;
         mem[864] = -13'h0003;
         mem[865] = -13'h00a5;
         mem[866] =  13'h0073;
         mem[867] =  13'h00bb;
         mem[868] =  13'h00a2;
         mem[869] =  13'h00ce;
         mem[870] = -13'h0046;
         mem[871] =  13'h0148;
         mem[872] =  13'h0190;
         mem[873] = -13'h003f;
         mem[874] = -13'h003e;
         mem[875] = -13'h0043;
         mem[876] = -13'h006b;
         mem[877] =  13'h0024;
         mem[878] = -13'h006e;
         mem[879] =  13'h001f;
         mem[880] = -13'h0041;
         mem[881] =  13'h0055;
         mem[882] =  13'h015e;
         mem[883] =  13'h0061;
         mem[884] = -13'h00a0;
         mem[885] = -13'h013f;
         mem[886] = -13'h0045;
         mem[887] =  13'h01e6;
         mem[888] =  13'h027f;
         mem[889] = -13'h00bc;
         mem[890] = -13'h002a;
         mem[891] =  13'h0188;
         mem[892] =  13'h0038;
         mem[893] =  13'h0009;
         mem[894] =  13'h0088;
         mem[895] = -13'h0088;
         mem[896] =  13'h000b;
         mem[897] = -13'h010d;
         mem[898] =  13'h0008;
         mem[899] =  13'h005b;
         mem[900] = -13'h00eb;
         mem[901] =  13'h001b;
         mem[902] =  13'h0032;
         mem[903] = -13'h0021;
         mem[904] =  13'h0096;
         mem[905] = -13'h066f;
         mem[906] = -13'h005a;
         mem[907] = -13'h0035;
         mem[908] = -13'h0034;
         mem[909] =  13'h0058;
         mem[910] =  13'h0030;
         mem[911] = -13'h0050;
         mem[912] =  13'h0107;
         mem[913] =  13'h01be;
         mem[914] = -13'h008b;
         mem[915] = -13'h000f;
         mem[916] = -13'h002c;
         mem[917] = -13'h002f;
         mem[918] =  13'h006a;
         mem[919] =  13'h0011;
         mem[920] = -13'h00c3;
         mem[921] =  13'h0001;
         mem[922] =  13'h01d8;
         mem[923] =  13'h0041;
         mem[924] =  13'h00e7;
         mem[925] = -13'h002b;
         mem[926] =  13'h01fc;
         mem[927] = -13'h0016;
         mem[928] =  13'h0030;
         mem[929] = -13'h00b0;
         mem[930] = -13'h0087;
         mem[931] = -13'h0057;
         mem[932] = -13'h0032;
         mem[933] = -13'h0045;
         mem[934] = -13'h000a;
         mem[935] = -13'h00b8;
         mem[936] =  13'h009f;
         mem[937] =  13'h001b;
         mem[938] = -13'h0043;
         mem[939] =  13'h0019;
         mem[940] =  13'h00bb;
         mem[941] =  13'h0010;
         mem[942] =  13'h0000;
         mem[943] =  13'h001d;
         mem[944] = -13'h00cc;
         mem[945] = -13'h0066;
         mem[946] =  13'h007e;
         mem[947] =  13'h00bd;
         mem[948] = -13'h000d;
         mem[949] = -13'h0063;
         mem[950] =  13'h0031;
         mem[951] =  13'h0035;
         mem[952] =  13'h00f2;
         mem[953] = -13'h00a8;
         mem[954] = -13'h0158;
         mem[955] =  13'h00b6;
         mem[956] =  13'h0064;
         mem[957] = -13'h0011;
         mem[958] =  13'h0064;
         mem[959] = -13'h015c;
         mem[960] =  13'h0059;
         mem[961] = -13'h0044;
         mem[962] =  13'h0085;
         mem[963] =  13'h000a;
         mem[964] =  13'h00e2;
         mem[965] = -13'h01b3;
         mem[966] = -13'h0020;
         mem[967] =  13'h0135;
         mem[968] = -13'h017c;
         mem[969] =  13'h00ca;
         mem[970] = -13'h0030;
         mem[971] =  13'h015f;
         mem[972] =  13'h014b;
         mem[973] = -13'h008a;
         mem[974] =  13'h003f;
         mem[975] =  13'h00e0;
         mem[976] =  13'h0057;
         mem[977] =  13'h0020;
         mem[978] = -13'h0099;
         mem[979] =  13'h028c;
         mem[980] = -13'h011a;
         mem[981] = -13'h008a;
         mem[982] = -13'h0103;
         mem[983] =  13'h001e;
         mem[984] = -13'h0027;
         mem[985] = -13'h0217;
         mem[986] =  13'h00eb;
         mem[987] = -13'h001d;
         mem[988] =  13'h007f;
         mem[989] =  13'h0092;
         mem[990] = -13'h0081;
         mem[991] = -13'h004f;
         mem[992] = -13'h001d;
         mem[993] =  13'h0021;
         mem[994] = -13'h00b2;
         mem[995] =  13'h006c;
         mem[996] =  13'h0083;
         mem[997] = -13'h0127;
         mem[998] =  13'h0080;
         mem[999] = -13'h0001;
         mem[1000] =  13'h000b;
         mem[1001] =  13'h0086;
         mem[1002] = -13'h003b;
         mem[1003] =  13'h009b;
         mem[1004] =  13'h000b;
         mem[1005] = -13'h00aa;
         mem[1006] = -13'h0065;
         mem[1007] =  13'h0029;
         mem[1008] = -13'h0055;
         mem[1009] =  13'h005b;
         mem[1010] = -13'h0098;
         mem[1011] = -13'h002b;
         mem[1012] =  13'h00e3;
         mem[1013] =  13'h0058;
         mem[1014] =  13'h0000;
         mem[1015] =  13'h003b;
         mem[1016] =  13'h01b9;
         mem[1017] =  13'h0093;
         mem[1018] = -13'h0010;
         mem[1019] =  13'h0055;
         mem[1020] = -13'h007a;
         mem[1021] =  13'h006a;
         mem[1022] =  13'h002b;
         mem[1023] =  13'h0023;
         mem[1024] =  13'h0057;
         mem[1025] =  13'h0131;
         mem[1026] =  13'h0013;
         mem[1027] =  13'h0007;
         mem[1028] =  13'h0004;
         mem[1029] =  13'h0073;
         mem[1030] = -13'h0085;
         mem[1031] =  13'h005c;
         mem[1032] = -13'h0058;
         mem[1033] =  13'h001f;
         mem[1034] =  13'h003b;
         mem[1035] =  13'h0072;
         mem[1036] =  13'h0017;
         mem[1037] = -13'h0028;
         mem[1038] = -13'h0010;
         mem[1039] = -13'h005c;
         mem[1040] = -13'h00a2;
         mem[1041] = -13'h0047;
         mem[1042] =  13'h0024;
         mem[1043] = -13'h0020;
         mem[1044] =  13'h006e;
         mem[1045] = -13'h0054;
         mem[1046] = -13'h0126;
         mem[1047] = -13'h006e;
         mem[1048] = -13'h00c2;
         mem[1049] = -13'h01be;
         mem[1050] =  13'h0037;
         mem[1051] = -13'h001b;
         mem[1052] = -13'h0010;
         mem[1053] = -13'h009a;
         mem[1054] =  13'h0023;
         mem[1055] = -13'h0083;
         mem[1056] =  13'h00ef;
         mem[1057] = -13'h00a7;
         mem[1058] = -13'h0051;
         mem[1059] = -13'h0012;
         mem[1060] =  13'h0044;
         mem[1061] =  13'h0026;
         mem[1062] = -13'h0050;
         mem[1063] =  13'h002c;
         mem[1064] =  13'h009b;
         mem[1065] =  13'h0043;
         mem[1066] = -13'h0051;
         mem[1067] =  13'h002d;
         mem[1068] =  13'h0015;
         mem[1069] = -13'h002d;
         mem[1070] = -13'h002b;
         mem[1071] =  13'h01af;
         mem[1072] =  13'h00e0;
         mem[1073] =  13'h0048;
         mem[1074] = -13'h007f;
         mem[1075] = -13'h00ea;
         mem[1076] = -13'h002e;
         mem[1077] =  13'h007d;
         mem[1078] =  13'h0007;
         mem[1079] =  13'h002e;
         mem[1080] =  13'h014d;
         mem[1081] =  13'h00db;
         mem[1082] = -13'h0062;
         mem[1083] =  13'h001b;
         mem[1084] = -13'h0084;
         mem[1085] =  13'h009b;
         mem[1086] =  13'h003f;
         mem[1087] = -13'h00b5;
         mem[1088] = -13'h005e;
         mem[1089] =  13'h004f;
         mem[1090] =  13'h01a9;
         mem[1091] = -13'h004d;
         mem[1092] =  13'h009e;
         mem[1093] =  13'h005d;
         mem[1094] = -13'h0080;
         mem[1095] =  13'h0027;
         mem[1096] = -13'h00c9;
         mem[1097] = -13'h00a1;
         mem[1098] =  13'h00c4;
         mem[1099] =  13'h00d2;
         mem[1100] =  13'h003a;
         mem[1101] = -13'h0177;
         mem[1102] =  13'h001a;
         mem[1103] =  13'h0092;
         mem[1104] =  13'h00cf;
         mem[1105] = -13'h003b;
         mem[1106] = -13'h009e;
         mem[1107] = -13'h00a5;
         mem[1108] =  13'h0061;
         mem[1109] =  13'h0023;
         mem[1110] = -13'h0220;
         mem[1111] =  13'h0028;
         mem[1112] =  13'h0014;
         mem[1113] = -13'h00fa;
         mem[1114] = -13'h0001;
         mem[1115] =  13'h000d;
         mem[1116] =  13'h0056;
         mem[1117] =  13'h001e;
         mem[1118] =  13'h0065;
         mem[1119] = -13'h0091;
         mem[1120] =  13'h0051;
         mem[1121] =  13'h003d;
         mem[1122] = -13'h005e;
         mem[1123] = -13'h004c;
         mem[1124] =  13'h0736;
         mem[1125] =  13'h0030;
         mem[1126] = -13'h0065;
         mem[1127] = -13'h00b7;
         mem[1128] = -13'h003b;
         mem[1129] = -13'h0064;
         mem[1130] =  13'h005e;
         mem[1131] = -13'h0066;
         mem[1132] =  13'h0004;
         mem[1133] =  13'h003f;
         mem[1134] = -13'h006d;
         mem[1135] =  13'h0005;
         mem[1136] = -13'h0002;
         mem[1137] = -13'h0082;
         mem[1138] = -13'h0014;
         mem[1139] =  13'h007f;
         mem[1140] = -13'h0089;
         mem[1141] =  13'h0031;
         mem[1142] = -13'h008e;
         mem[1143] =  13'h0028;
         mem[1144] =  13'h00f4;
         mem[1145] = -13'h010b;
         mem[1146] = -13'h017c;
         mem[1147] = -13'h00a8;
         mem[1148] =  13'h0057;
         mem[1149] = -13'h0068;
         mem[1150] = -13'h00a8;
         mem[1151] = -13'h0048;
         mem[1152] =  13'h0024;
         mem[1153] = -13'h002f;
         mem[1154] = -13'h001e;
         mem[1155] =  13'h0003;
         mem[1156] = -13'h007d;
         mem[1157] = -13'h004d;
         mem[1158] = -13'h0021;
         mem[1159] = -13'h008e;
         mem[1160] =  13'h004d;
         mem[1161] = -13'h004d;
         mem[1162] = -13'h016c;
         mem[1163] =  13'h001c;
         mem[1164] = -13'h0073;
         mem[1165] = -13'h0001;
         mem[1166] = -13'h01bb;
         mem[1167] =  13'h0041;
         mem[1168] =  13'h0023;
         mem[1169] = -13'h0067;
         mem[1170] = -13'h0037;
         mem[1171] = -13'h001f;
         mem[1172] =  13'h0125;
         mem[1173] = -13'h0037;
         mem[1174] =  13'h000c;
         mem[1175] = -13'h00d0;
         mem[1176] = -13'h0024;
         mem[1177] =  13'h036d;
         mem[1178] =  13'h0039;
         mem[1179] =  13'h00ae;
         mem[1180] =  13'h0051;
         mem[1181] = -13'h0089;
         mem[1182] =  13'h0104;
         mem[1183] =  13'h0059;
         mem[1184] = -13'h0141;
         mem[1185] =  13'h003a;
         mem[1186] = -13'h0113;
         mem[1187] =  13'h0216;
         mem[1188] = -13'h00bd;
         mem[1189] = -13'h007a;
         mem[1190] = -13'h0001;
         mem[1191] = -13'h005b;
         mem[1192] = -13'h0006;
         mem[1193] =  13'h0031;
         mem[1194] =  13'h0063;
         mem[1195] = -13'h00c1;
         mem[1196] = -13'h0065;
         mem[1197] =  13'h0059;
         mem[1198] =  13'h0302;
         mem[1199] = -13'h013e;
         mem[1200] = -13'h00c7;
         mem[1201] = -13'h0046;
         mem[1202] = -13'h000b;
         mem[1203] = -13'h0194;
         mem[1204] = -13'h0059;
         mem[1205] =  13'h00fa;
         mem[1206] = -13'h0064;
         mem[1207] =  13'h008a;
         mem[1208] =  13'h009c;
         mem[1209] = -13'h0052;
         mem[1210] =  13'h0065;
         mem[1211] = -13'h0063;
         mem[1212] = -13'h006c;
         mem[1213] = -13'h000e;
         mem[1214] =  13'h01b6;
         mem[1215] =  13'h00b8;
         mem[1216] =  13'h00b5;
         mem[1217] =  13'h0004;
         mem[1218] =  13'h0124;
         mem[1219] =  13'h0092;
         mem[1220] = -13'h0055;
         mem[1221] =  13'h06cd;
         mem[1222] =  13'h002e;
         mem[1223] = -13'h003e;
         mem[1224] = -13'h003e;
         mem[1225] = -13'h004d;
         mem[1226] = -13'h000d;
         mem[1227] =  13'h017d;
         mem[1228] = -13'h0033;
         mem[1229] = -13'h006e;
         mem[1230] = -13'h0060;
         mem[1231] = -13'h003a;
         mem[1232] =  13'h0073;
         mem[1233] =  13'h00d0;
         mem[1234] =  13'h002f;
         mem[1235] = -13'h003c;
         mem[1236] =  13'h03a7;
         mem[1237] =  13'h01c6;
         mem[1238] =  13'h000d;
         mem[1239] =  13'h015d;
         mem[1240] =  13'h005a;
         mem[1241] = -13'h0040;
         mem[1242] =  13'h054c;
         mem[1243] =  13'h0024;
         mem[1244] =  13'h00bc;
         mem[1245] = -13'h009a;
         mem[1246] = -13'h014f;
         mem[1247] =  13'h037b;
         mem[1248] =  13'h003c;
         mem[1249] =  13'h00d6;
         mem[1250] =  13'h0025;
         mem[1251] =  13'h0020;
         mem[1252] = -13'h006a;
         mem[1253] = -13'h000c;
         mem[1254] =  13'h00ea;
         mem[1255] = -13'h0019;
         mem[1256] = -13'h00a5;
         mem[1257] = -13'h0053;
         mem[1258] = -13'h0046;
         mem[1259] = -13'h0063;
         mem[1260] =  13'h00e8;
         mem[1261] =  13'h0001;
         mem[1262] =  13'h0028;
         mem[1263] = -13'h00d7;
         mem[1264] = -13'h0038;
         mem[1265] = -13'h007c;
         mem[1266] = -13'h04ce;
         mem[1267] = -13'h0093;
         mem[1268] = -13'h00e1;
         mem[1269] =  13'h008a;
         mem[1270] = -13'h0021;
         mem[1271] = -13'h0016;
         mem[1272] =  13'h000c;
         mem[1273] =  13'h00db;
         mem[1274] = -13'h0201;
         mem[1275] =  13'h017b;
         mem[1276] =  13'h009d;
         mem[1277] = -13'h0008;
         mem[1278] =  13'h0027;
         mem[1279] =  13'h0062;
         mem[1280] = -13'h0049;
         mem[1281] = -13'h002b;
         mem[1282] = -13'h001d;
         mem[1283] =  13'h0062;
         mem[1284] = -13'h004b;
         mem[1285] =  13'h0040;
         mem[1286] = -13'h00c7;
         mem[1287] =  13'h001b;
         mem[1288] =  13'h0028;
         mem[1289] =  13'h003c;
         mem[1290] =  13'h018d;
         mem[1291] =  13'h00c5;
         mem[1292] =  13'h0028;
         mem[1293] = -13'h00a3;
         mem[1294] =  13'h005d;
         mem[1295] =  13'h001b;
         mem[1296] =  13'h00f4;
         mem[1297] =  13'h001c;
         mem[1298] =  13'h0040;
         mem[1299] = -13'h00cb;
         mem[1300] =  13'h00d6;
         mem[1301] =  13'h005b;
         mem[1302] =  13'h00a8;
         mem[1303] = -13'h0058;
         mem[1304] = -13'h0153;
         mem[1305] =  13'h0022;
         mem[1306] =  13'h0143;
         mem[1307] = -13'h0171;
         mem[1308] = -13'h0077;
         mem[1309] =  13'h001c;
         mem[1310] = -13'h0021;
         mem[1311] =  13'h0050;
         mem[1312] = -13'h003c;
         mem[1313] =  13'h0067;
         mem[1314] = -13'h0040;
         mem[1315] =  13'h0078;
         mem[1316] = -13'h0022;
         mem[1317] =  13'h0064;
         mem[1318] = -13'h008a;
         mem[1319] = -13'h0008;
         mem[1320] =  13'h007c;
         mem[1321] =  13'h0010;
         mem[1322] =  13'h0071;
         mem[1323] =  13'h0020;
         mem[1324] =  13'h00b4;
         mem[1325] = -13'h0084;
         mem[1326] =  13'h0055;
         mem[1327] =  13'h0067;
         mem[1328] =  13'h001a;
         mem[1329] = -13'h00ef;
         mem[1330] =  13'h0082;
         mem[1331] = -13'h007c;
         mem[1332] =  13'h003d;
         mem[1333] = -13'h00c8;
         mem[1334] =  13'h0154;
         mem[1335] =  13'h0061;
         mem[1336] =  13'h0043;
         mem[1337] = -13'h0030;
         mem[1338] =  13'h0000;
         mem[1339] =  13'h004e;
         mem[1340] = -13'h0029;
         mem[1341] = -13'h0039;
         mem[1342] = -13'h01a6;
         mem[1343] = -13'h0187;
         mem[1344] = -13'h00a9;
         mem[1345] =  13'h0009;
         mem[1346] =  13'h01b7;
         mem[1347] =  13'h000d;
         mem[1348] =  13'h0077;
         mem[1349] =  13'h002e;
         mem[1350] = -13'h0031;
         mem[1351] = -13'h0034;
         mem[1352] =  13'h0064;
         mem[1353] =  13'h00bc;
         mem[1354] = -13'h006f;
         mem[1355] =  13'h00a4;
         mem[1356] =  13'h005e;
         mem[1357] = -13'h0061;
         mem[1358] =  13'h013d;
         mem[1359] = -13'h0036;
         mem[1360] = -13'h0058;
         mem[1361] = -13'h0124;
         mem[1362] = -13'h0016;
         mem[1363] =  13'h006d;
         mem[1364] = -13'h00a1;
         mem[1365] =  13'h006a;
         mem[1366] =  13'h00c8;
         mem[1367] =  13'h0097;
         mem[1368] =  13'h0143;
         mem[1369] =  13'h0076;
         mem[1370] =  13'h0019;
         mem[1371] = -13'h010d;
         mem[1372] = -13'h011a;
         mem[1373] = -13'h01dd;
         mem[1374] = -13'h0005;
         mem[1375] = -13'h00b6;
         mem[1376] =  13'h00d1;
         mem[1377] = -13'h0081;
         mem[1378] =  13'h0056;
         mem[1379] = -13'h0236;
         mem[1380] =  13'h00d5;
         mem[1381] =  13'h006a;
         mem[1382] = -13'h0031;
         mem[1383] = -13'h0063;
         mem[1384] = -13'h0067;
         mem[1385] =  13'h0033;
         mem[1386] =  13'h00ea;
         mem[1387] =  13'h0044;
         mem[1388] = -13'h005d;
         mem[1389] =  13'h0000;
         mem[1390] = -13'h001f;
         mem[1391] =  13'h0181;
         mem[1392] = -13'h00ff;
         mem[1393] =  13'h0047;
         mem[1394] = -13'h005a;
         mem[1395] = -13'h002a;
         mem[1396] = -13'h0026;
         mem[1397] = -13'h0076;
         mem[1398] = -13'h0056;
         mem[1399] = -13'h0097;
         mem[1400] =  13'h002b;
         mem[1401] =  13'h029e;
         mem[1402] =  13'h0184;
         mem[1403] =  13'h0090;
         mem[1404] =  13'h0034;
         mem[1405] =  13'h0239;
         mem[1406] =  13'h0030;
         mem[1407] = -13'h0028;
         mem[1408] = -13'h0018;
         mem[1409] = -13'h0005;
         mem[1410] =  13'h0084;
         mem[1411] = -13'h0039;
         mem[1412] =  13'h0004;
         mem[1413] =  13'h0000;
         mem[1414] = -13'h0001;
         mem[1415] =  13'h0010;
         mem[1416] =  13'h003a;
         mem[1417] = -13'h00e2;
         mem[1418] =  13'h017f;
         mem[1419] =  13'h006d;
         mem[1420] =  13'h000f;
         mem[1421] = -13'h0082;
         mem[1422] = -13'h005c;
         mem[1423] =  13'h0067;
         mem[1424] = -13'h007f;
         mem[1425] = -13'h006c;
         mem[1426] = -13'h0038;
         mem[1427] = -13'h0101;
         mem[1428] = -13'h00b7;
         mem[1429] = -13'h0053;
         mem[1430] = -13'h0020;
         mem[1431] =  13'h0023;
         mem[1432] = -13'h006f;
         mem[1433] = -13'h0043;
         mem[1434] = -13'h0038;
         mem[1435] =  13'h0077;
         mem[1436] =  13'h0099;
         mem[1437] = -13'h0066;
         mem[1438] = -13'h0105;
         mem[1439] = -13'h0026;
         mem[1440] = -13'h0003;
         mem[1441] = -13'h0059;
         mem[1442] = -13'h0049;
         mem[1443] = -13'h0065;
         mem[1444] =  13'h0283;
         mem[1445] =  13'h011a;
         mem[1446] = -13'h002d;
         mem[1447] = -13'h0038;
         mem[1448] = -13'h007e;
         mem[1449] =  13'h0057;
         mem[1450] =  13'h017d;
         mem[1451] =  13'h0079;
         mem[1452] =  13'h0000;
         mem[1453] = -13'h00ac;
         mem[1454] = -13'h005c;
         mem[1455] = -13'h0034;
         mem[1456] =  13'h0072;
         mem[1457] = -13'h0071;
         mem[1458] = -13'h0019;
         mem[1459] = -13'h0053;
         mem[1460] = -13'h0032;
         mem[1461] = -13'h00a5;
         mem[1462] =  13'h0079;
         mem[1463] =  13'h001c;
         mem[1464] =  13'h0042;
         mem[1465] =  13'h00cd;
         mem[1466] =  13'h0008;
         mem[1467] =  13'h0066;
         mem[1468] = -13'h0040;
         mem[1469] =  13'h0098;
         mem[1470] = -13'h0144;
         mem[1471] = -13'h0046;
         mem[1472] =  13'h0086;
         mem[1473] = -13'h01e1;
         mem[1474] =  13'h01ed;
         mem[1475] =  13'h0011;
         mem[1476] = -13'h0129;
         mem[1477] =  13'h02d5;
         mem[1478] =  13'h0022;
         mem[1479] = -13'h0035;
         mem[1480] =  13'h004d;
         mem[1481] =  13'h0057;
         mem[1482] =  13'h0103;
         mem[1483] = -13'h0084;
         mem[1484] = -13'h0060;
         mem[1485] =  13'h004c;
         mem[1486] =  13'h007f;
         mem[1487] = -13'h002d;
         mem[1488] = -13'h0034;
         mem[1489] = -13'h0034;
         mem[1490] =  13'h0119;
         mem[1491] =  13'h0015;
         mem[1492] = -13'h009e;
         mem[1493] =  13'h0019;
         mem[1494] =  13'h02cd;
         mem[1495] =  13'h01dc;
         mem[1496] = -13'h005e;
         mem[1497] = -13'h00d2;
         mem[1498] =  13'h0398;
         mem[1499] =  13'h0026;
         mem[1500] = -13'h01e5;
         mem[1501] =  13'h009a;
         mem[1502] =  13'h005a;
         mem[1503] = -13'h0094;
         mem[1504] = -13'h021c;
         mem[1505] = -13'h00aa;
         mem[1506] = -13'h0087;
         mem[1507] =  13'h0040;
         mem[1508] = -13'h00a1;
         mem[1509] = -13'h0115;
         mem[1510] = -13'h006d;
         mem[1511] =  13'h00a3;
         mem[1512] =  13'h019c;
         mem[1513] = -13'h014b;
         mem[1514] = -13'h0057;
         mem[1515] = -13'h002b;
         mem[1516] =  13'h0003;
         mem[1517] =  13'h000e;
         mem[1518] =  13'h004d;
         mem[1519] = -13'h0068;
         mem[1520] = -13'h0010;
         mem[1521] = -13'h0003;
         mem[1522] = -13'h00ca;
         mem[1523] =  13'h002f;
         mem[1524] =  13'h008d;
         mem[1525] = -13'h0021;
         mem[1526] = -13'h005b;
         mem[1527] = -13'h007e;
         mem[1528] =  13'h00b3;
         mem[1529] =  13'h00b0;
         mem[1530] =  13'h006f;
         mem[1531] =  13'h0026;
         mem[1532] =  13'h0182;
         mem[1533] =  13'h02b9;
         mem[1534] = -13'h00c1;
         mem[1535] =  13'h01ca;
         mem[1536] = -13'h003a;
         mem[1537] =  13'h008b;
         mem[1538] =  13'h0058;
         mem[1539] =  13'h0059;
         mem[1540] =  13'h0151;
         mem[1541] =  13'h015a;
         mem[1542] = -13'h00e1;
         mem[1543] = -13'h0109;
         mem[1544] = -13'h005d;
         mem[1545] =  13'h00e0;
         mem[1546] =  13'h0000;
         mem[1547] =  13'h0192;
         mem[1548] = -13'h001d;
         mem[1549] =  13'h00cd;
         mem[1550] = -13'h0017;
         mem[1551] =  13'h0039;
         mem[1552] =  13'h0057;
         mem[1553] = -13'h0077;
         mem[1554] =  13'h0001;
         mem[1555] =  13'h0007;
         mem[1556] =  13'h0023;
         mem[1557] =  13'h0104;
         mem[1558] = -13'h0072;
         mem[1559] =  13'h00c8;
         mem[1560] = -13'h0078;
         mem[1561] =  13'h01fc;
         mem[1562] =  13'h0020;
         mem[1563] =  13'h007c;
         mem[1564] =  13'h0067;
         mem[1565] =  13'h0029;
         mem[1566] = -13'h0044;
         mem[1567] = -13'h000b;
         mem[1568] =  13'h00ad;
         mem[1569] = -13'h00c6;
         mem[1570] =  13'h0076;
         mem[1571] = -13'h00a4;
         mem[1572] = -13'h00a8;
         mem[1573] =  13'h0030;
         mem[1574] = -13'h0057;
         mem[1575] = -13'h0061;
         mem[1576] =  13'h0049;
         mem[1577] = -13'h00b2;
         mem[1578] = -13'h0025;
         mem[1579] =  13'h00c2;
         mem[1580] = -13'h003a;
         mem[1581] =  13'h000f;
         mem[1582] =  13'h000e;
         mem[1583] = -13'h0077;
         mem[1584] = -13'h001a;
         mem[1585] = -13'h007b;
         mem[1586] =  13'h0020;
         mem[1587] =  13'h0024;
         mem[1588] =  13'h0189;
         mem[1589] = -13'h0086;
         mem[1590] = -13'h0036;
         mem[1591] =  13'h003e;
         mem[1592] =  13'h0031;
         mem[1593] = -13'h0138;
         mem[1594] = -13'h0031;
         mem[1595] =  13'h0059;
         mem[1596] = -13'h000b;
         mem[1597] = -13'h00c7;
         mem[1598] = -13'h002a;
         mem[1599] = -13'h001b;
         mem[1600] =  13'h0023;
         mem[1601] =  13'h0051;
         mem[1602] =  13'h005a;
         mem[1603] = -13'h00d5;
         mem[1604] =  13'h0050;
         mem[1605] =  13'h005e;
         mem[1606] = -13'h003d;
         mem[1607] = -13'h00cc;
         mem[1608] = -13'h011b;
         mem[1609] =  13'h0013;
         mem[1610] = -13'h008a;
         mem[1611] = -13'h0042;
         mem[1612] = -13'h00cd;
         mem[1613] =  13'h00e9;
         mem[1614] =  13'h00a7;
         mem[1615] = -13'h000c;
         mem[1616] = -13'h0085;
         mem[1617] =  13'h0193;
         mem[1618] = -13'h009c;
         mem[1619] = -13'h00bc;
         mem[1620] = -13'h01e9;
         mem[1621] = -13'h01ed;
         mem[1622] =  13'h0121;
         mem[1623] =  13'h0022;
         mem[1624] =  13'h005d;
         mem[1625] =  13'h0002;
         mem[1626] =  13'h008d;
         mem[1627] = -13'h0012;
         mem[1628] =  13'h0060;
         mem[1629] =  13'h0034;
         mem[1630] = -13'h002e;
         mem[1631] = -13'h00aa;
         mem[1632] = -13'h017e;
         mem[1633] = -13'h006f;
         mem[1634] = -13'h0059;
         mem[1635] = -13'h0027;
         mem[1636] =  13'h011c;
         mem[1637] =  13'h007f;
         mem[1638] = -13'h00cb;
         mem[1639] = -13'h0053;
         mem[1640] = -13'h003e;
         mem[1641] = -13'h00cf;
         mem[1642] = -13'h0054;
         mem[1643] = -13'h007e;
         mem[1644] = -13'h0012;
         mem[1645] = -13'h00bb;
         mem[1646] =  13'h0044;
         mem[1647] =  13'h000d;
         mem[1648] =  13'h0064;
         mem[1649] = -13'h0146;
         mem[1650] =  13'h00b6;
         mem[1651] = -13'h0201;
         mem[1652] =  13'h0049;
         mem[1653] =  13'h004e;
         mem[1654] =  13'h00a3;
         mem[1655] =  13'h0037;
         mem[1656] =  13'h0042;
         mem[1657] =  13'h002d;
         mem[1658] =  13'h00a0;
         mem[1659] = -13'h0027;
         mem[1660] =  13'h0072;
         mem[1661] = -13'h0060;
         mem[1662] =  13'h006e;
         mem[1663] =  13'h0001;
         mem[1664] = -13'h00a8;
         mem[1665] =  13'h001b;
         mem[1666] =  13'h00c4;
         mem[1667] = -13'h000c;
         mem[1668] = -13'h0023;
         mem[1669] = -13'h001e;
         mem[1670] = -13'h0007;
         mem[1671] = -13'h0161;
         mem[1672] =  13'h00bf;
         mem[1673] =  13'h0000;
         mem[1674] = -13'h0042;
         mem[1675] =  13'h00bb;
         mem[1676] = -13'h0070;
         mem[1677] = -13'h0071;
         mem[1678] =  13'h001f;
         mem[1679] = -13'h0002;
         mem[1680] =  13'h01c4;
         mem[1681] =  13'h0119;
         mem[1682] =  13'h0007;
         mem[1683] =  13'h0313;
         mem[1684] =  13'h0284;
         mem[1685] = -13'h00ca;
         mem[1686] =  13'h00d4;
         mem[1687] =  13'h00cc;
         mem[1688] = -13'h00ae;
         mem[1689] = -13'h0099;
         mem[1690] = -13'h0098;
         mem[1691] =  13'h0039;
         mem[1692] = -13'h0001;
         mem[1693] =  13'h0083;
         mem[1694] = -13'h0011;
         mem[1695] =  13'h0028;
         mem[1696] =  13'h017e;
         mem[1697] =  13'h0046;
         mem[1698] =  13'h0022;
         mem[1699] = -13'h0039;
         mem[1700] = -13'h001f;
         mem[1701] =  13'h0072;
         mem[1702] = -13'h004d;
         mem[1703] = -13'h004c;
         mem[1704] = -13'h0095;
         mem[1705] =  13'h0084;
         mem[1706] =  13'h00f4;
         mem[1707] =  13'h0028;
         mem[1708] = -13'h0090;
         mem[1709] =  13'h000b;
         mem[1710] =  13'h0021;
         mem[1711] =  13'h016c;
         mem[1712] = -13'h007b;
         mem[1713] = -13'h0059;
         mem[1714] =  13'h009a;
         mem[1715] =  13'h000b;
         mem[1716] = -13'h002b;
         mem[1717] =  13'h0213;
         mem[1718] = -13'h0048;
         mem[1719] = -13'h013b;
         mem[1720] = -13'h004e;
         mem[1721] = -13'h00d1;
         mem[1722] =  13'h0008;
         mem[1723] =  13'h0068;
         mem[1724] = -13'h0061;
         mem[1725] = -13'h001a;
         mem[1726] = -13'h009a;
         mem[1727] =  13'h0376;
         mem[1728] = -13'h0036;
         mem[1729] =  13'h0123;
         mem[1730] =  13'h00e5;
         mem[1731] =  13'h00a5;
         mem[1732] =  13'h0102;
         mem[1733] =  13'h002a;
         mem[1734] =  13'h0100;
         mem[1735] = -13'h00a1;
         mem[1736] = -13'h0016;
         mem[1737] =  13'h01b9;
         mem[1738] =  13'h0045;
         mem[1739] =  13'h007f;
         mem[1740] = -13'h005e;
         mem[1741] = -13'h002d;
         mem[1742] = -13'h0013;
         mem[1743] = -13'h0047;
         mem[1744] =  13'h004d;
         mem[1745] =  13'h001d;
         mem[1746] =  13'h004d;
         mem[1747] =  13'h007f;
         mem[1748] =  13'h0055;
         mem[1749] =  13'h002e;
         mem[1750] = -13'h00e9;
         mem[1751] =  13'h0127;
         mem[1752] = -13'h0051;
         mem[1753] = -13'h0044;
         mem[1754] = -13'h00a3;
         mem[1755] =  13'h006e;
         mem[1756] = -13'h0010;
         mem[1757] =  13'h005d;
         mem[1758] = -13'h011a;
         mem[1759] =  13'h00b0;
         mem[1760] =  13'h0023;
         mem[1761] =  13'h003b;
         mem[1762] = -13'h002f;
         mem[1763] = -13'h01c1;
         mem[1764] =  13'h00b9;
         mem[1765] = -13'h006e;
         mem[1766] =  13'h0049;
         mem[1767] =  13'h00ce;
         mem[1768] = -13'h007a;
         mem[1769] =  13'h009b;
         mem[1770] =  13'h02f8;
         mem[1771] = -13'h0010;
         mem[1772] =  13'h0029;
         mem[1773] = -13'h002f;
         mem[1774] = -13'h001a;
         mem[1775] =  13'h002b;
         mem[1776] = -13'h0053;
         mem[1777] =  13'h0009;
         mem[1778] = -13'h0006;
         mem[1779] =  13'h0023;
         mem[1780] = -13'h0063;
         mem[1781] =  13'h0130;
         mem[1782] =  13'h0045;
         mem[1783] = -13'h0064;
         mem[1784] =  13'h007b;
         mem[1785] =  13'h0031;
         mem[1786] =  13'h0163;
         mem[1787] = -13'h00ad;
         mem[1788] = -13'h000a;
         mem[1789] = -13'h00e8;
         mem[1790] =  13'h0060;
         mem[1791] = -13'h0055;
         mem[1792] =  13'h001d;
         mem[1793] =  13'h0577;
         mem[1794] =  13'h0019;
         mem[1795] =  13'h0085;
         mem[1796] =  13'h0000;
         mem[1797] =  13'h0002;
         mem[1798] =  13'h00df;
         mem[1799] = -13'h0029;
         mem[1800] = -13'h004d;
         mem[1801] = -13'h0015;
         mem[1802] = -13'h002c;
         mem[1803] = -13'h00cc;
         mem[1804] =  13'h0031;
         mem[1805] = -13'h0009;
         mem[1806] =  13'h000c;
         mem[1807] =  13'h0010;
         mem[1808] = -13'h001e;
         mem[1809] =  13'h00d4;
         mem[1810] =  13'h004b;
         mem[1811] =  13'h02cc;
         mem[1812] =  13'h00dd;
         mem[1813] = -13'h0520;
         mem[1814] = -13'h006e;
         mem[1815] =  13'h013d;
         mem[1816] =  13'h0061;
         mem[1817] =  13'h002f;
         mem[1818] =  13'h0085;
         mem[1819] = -13'h00b5;
         mem[1820] = -13'h00ef;
         mem[1821] =  13'h004f;
         mem[1822] = -13'h00b7;
         mem[1823] = -13'h00f7;
         mem[1824] =  13'h002f;
         mem[1825] =  13'h0072;
         mem[1826] =  13'h010b;
         mem[1827] =  13'h0027;
         mem[1828] =  13'h000a;
         mem[1829] =  13'h0082;
         mem[1830] =  13'h0087;
         mem[1831] =  13'h00c2;
         mem[1832] = -13'h0050;
         mem[1833] = -13'h00e0;
         mem[1834] = -13'h005c;
         mem[1835] =  13'h01b6;
         mem[1836] = -13'h0095;
         mem[1837] =  13'h0039;
         mem[1838] =  13'h0055;
         mem[1839] =  13'h00c9;
         mem[1840] =  13'h0094;
         mem[1841] =  13'h00a8;
         mem[1842] =  13'h0040;
         mem[1843] = -13'h0042;
         mem[1844] = -13'h000c;
         mem[1845] = -13'h0234;
         mem[1846] = -13'h0027;
         mem[1847] = -13'h0065;
         mem[1848] = -13'h023b;
         mem[1849] = -13'h0150;
         mem[1850] =  13'h000f;
         mem[1851] = -13'h001b;
         mem[1852] = -13'h0041;
         mem[1853] = -13'h00d0;
         mem[1854] =  13'h0044;
         mem[1855] =  13'h0041;
         mem[1856] =  13'h000e;
         mem[1857] = -13'h0160;
         mem[1858] =  13'h0087;
         mem[1859] = -13'h0010;
         mem[1860] = -13'h0062;
         mem[1861] =  13'h0023;
         mem[1862] = -13'h0071;
         mem[1863] = -13'h031c;
         mem[1864] = -13'h01bd;
         mem[1865] = -13'h004f;
         mem[1866] =  13'h000c;
         mem[1867] =  13'h00f2;
         mem[1868] = -13'h00de;
         mem[1869] = -13'h00a1;
         mem[1870] =  13'h0151;
         mem[1871] = -13'h001e;
         mem[1872] =  13'h001e;
         mem[1873] =  13'h001c;
         mem[1874] = -13'h003f;
         mem[1875] = -13'h000b;
         mem[1876] = -13'h0121;
         mem[1877] = -13'h002f;
         mem[1878] =  13'h0002;
         mem[1879] = -13'h0097;
         mem[1880] = -13'h0085;
         mem[1881] = -13'h0132;
         mem[1882] =  13'h00a9;
         mem[1883] = -13'h0076;
         mem[1884] =  13'h00bd;
         mem[1885] =  13'h0411;
         mem[1886] =  13'h0009;
         mem[1887] = -13'h0153;
         mem[1888] = -13'h002e;
         mem[1889] = -13'h0210;
         mem[1890] =  13'h009d;
         mem[1891] =  13'h01a1;
         mem[1892] = -13'h004e;
         mem[1893] = -13'h00f8;
         mem[1894] =  13'h0065;
         mem[1895] =  13'h006d;
         mem[1896] =  13'h003d;
         mem[1897] =  13'h006b;
         mem[1898] = -13'h0099;
         mem[1899] = -13'h0015;
         mem[1900] =  13'h0048;
         mem[1901] = -13'h008b;
         mem[1902] = -13'h0041;
         mem[1903] =  13'h0050;
         mem[1904] = -13'h01a8;
         mem[1905] = -13'h004e;
         mem[1906] = -13'h0034;
         mem[1907] = -13'h0042;
         mem[1908] = -13'h020a;
         mem[1909] =  13'h004e;
         mem[1910] =  13'h0085;
         mem[1911] =  13'h0026;
         mem[1912] =  13'h0014;
         mem[1913] =  13'h00a9;
         mem[1914] = -13'h0138;
         mem[1915] = -13'h012a;
         mem[1916] =  13'h00f4;
         mem[1917] =  13'h0053;
         mem[1918] = -13'h0148;
         mem[1919] = -13'h0049;
         mem[1920] =  13'h002e;
         mem[1921] = -13'h0068;
         mem[1922] = -13'h0003;
         mem[1923] = -13'h003b;
         mem[1924] =  13'h0023;
         mem[1925] =  13'h00e0;
         mem[1926] = -13'h01bb;
         mem[1927] =  13'h005e;
         mem[1928] =  13'h000b;
         mem[1929] = -13'h0008;
         mem[1930] = -13'h005c;
         mem[1931] =  13'h0154;
         mem[1932] = -13'h001b;
         mem[1933] =  13'h0139;
         mem[1934] =  13'h0016;
         mem[1935] = -13'h002a;
         mem[1936] =  13'h0071;
         mem[1937] = -13'h005f;
         mem[1938] = -13'h00e3;
         mem[1939] = -13'h00a6;
         mem[1940] = -13'h001e;
         mem[1941] =  13'h0045;
         mem[1942] = -13'h0097;
         mem[1943] = -13'h0050;
         mem[1944] = -13'h0060;
         mem[1945] = -13'h00b1;
         mem[1946] = -13'h005a;
         mem[1947] =  13'h0043;
         mem[1948] = -13'h0086;
         mem[1949] =  13'h0124;
         mem[1950] =  13'h0003;
         mem[1951] = -13'h0022;
         mem[1952] = -13'h0046;
         mem[1953] = -13'h004c;
         mem[1954] = -13'h0025;
         mem[1955] =  13'h004b;
         mem[1956] = -13'h00ce;
         mem[1957] = -13'h0060;
         mem[1958] = -13'h006f;
         mem[1959] =  13'h001a;
         mem[1960] =  13'h005f;
         mem[1961] =  13'h0035;
         mem[1962] = -13'h001b;
         mem[1963] = -13'h005c;
         mem[1964] = -13'h0105;
         mem[1965] = -13'h00cc;
         mem[1966] =  13'h001b;
         mem[1967] = -13'h00e4;
         mem[1968] =  13'h051c;
         mem[1969] =  13'h014b;
         mem[1970] = -13'h003d;
         mem[1971] =  13'h00bf;
         mem[1972] =  13'h0018;
         mem[1973] = -13'h008c;
         mem[1974] = -13'h008f;
         mem[1975] =  13'h000c;
         mem[1976] = -13'h0039;
         mem[1977] = -13'h001b;
         mem[1978] = -13'h00d8;
         mem[1979] = -13'h0008;
         mem[1980] =  13'h004b;
         mem[1981] =  13'h0033;
         mem[1982] =  13'h0034;
         mem[1983] = -13'h0049;
         mem[1984] =  13'h0007;
         mem[1985] = -13'h003c;
         mem[1986] = -13'h003d;
         mem[1987] =  13'h003b;
         mem[1988] = -13'h002c;
         mem[1989] = -13'h0025;
         mem[1990] =  13'h0012;
         mem[1991] =  13'h0060;
         mem[1992] =  13'h0082;
         mem[1993] = -13'h004b;
         mem[1994] =  13'h0050;
         mem[1995] =  13'h0695;
         mem[1996] = -13'h00aa;
         mem[1997] = -13'h002a;
         mem[1998] =  13'h0032;
         mem[1999] = -13'h0023;
         mem[2000] =  13'h0042;
         mem[2001] = -13'h002a;
         mem[2002] = -13'h0032;
         mem[2003] = -13'h00ce;
         mem[2004] =  13'h00ca;
         mem[2005] = -13'h00a8;
         mem[2006] =  13'h0004;
         mem[2007] = -13'h00cd;
         mem[2008] = -13'h0023;
         mem[2009] = -13'h00cd;
         mem[2010] =  13'h01a2;
         mem[2011] = -13'h003a;
         mem[2012] =  13'h002a;
         mem[2013] = -13'h0030;
         mem[2014] =  13'h0127;
         mem[2015] = -13'h004d;
         mem[2016] = -13'h0013;
         mem[2017] = -13'h00ee;
         mem[2018] =  13'h0004;
         mem[2019] = -13'h00ca;
         mem[2020] = -13'h01e7;
         mem[2021] = -13'h004a;
         mem[2022] = -13'h0020;
         mem[2023] =  13'h00d4;
         mem[2024] =  13'h0111;
         mem[2025] = -13'h0038;
         mem[2026] = -13'h0048;
         mem[2027] = -13'h00ac;
         mem[2028] = -13'h0037;
         mem[2029] = -13'h002d;
         mem[2030] = -13'h01f7;
         mem[2031] =  13'h00c3;
         mem[2032] =  13'h0082;
         mem[2033] =  13'h0011;
         mem[2034] = -13'h00fb;
         mem[2035] = -13'h000b;
         mem[2036] = -13'h0118;
         mem[2037] =  13'h01a8;
         mem[2038] =  13'h0040;
         mem[2039] = -13'h0028;
         mem[2040] = -13'h0024;
         mem[2041] = -13'h0105;
         mem[2042] =  13'h009f;
         mem[2043] = -13'h00a3;
         mem[2044] =  13'h00ce;
         mem[2045] =  13'h00bd;
         mem[2046] =  13'h00fe;
         mem[2047] = -13'h0109;
         mem[2048] =  13'h0070;
         mem[2049] =  13'h0001;
         mem[2050] = -13'h0011;
         mem[2051] =  13'h00c1;
         mem[2052] =  13'h0033;
         mem[2053] =  13'h00bc;
         mem[2054] =  13'h032d;
         mem[2055] =  13'h0044;
         mem[2056] =  13'h0008;
         mem[2057] =  13'h005b;
         mem[2058] = -13'h0038;
         mem[2059] = -13'h001f;
         mem[2060] = -13'h0036;
         mem[2061] =  13'h00c8;
         mem[2062] =  13'h0053;
         mem[2063] = -13'h0044;
         mem[2064] = -13'h02b5;
         mem[2065] = -13'h01d0;
         mem[2066] = -13'h013e;
         mem[2067] = -13'h003f;
         mem[2068] = -13'h010e;
         mem[2069] =  13'h0022;
         mem[2070] =  13'h0091;
         mem[2071] = -13'h009f;
         mem[2072] = -13'h0028;
         mem[2073] = -13'h005e;
         mem[2074] =  13'h000c;
         mem[2075] =  13'h0035;
         mem[2076] =  13'h003c;
         mem[2077] = -13'h00f6;
         mem[2078] =  13'h00d4;
         mem[2079] =  13'h0065;
         mem[2080] = -13'h0031;
         mem[2081] = -13'h0194;
         mem[2082] =  13'h01e1;
         mem[2083] = -13'h004d;
         mem[2084] = -13'h0074;
         mem[2085] =  13'h0035;
         mem[2086] = -13'h01dd;
         mem[2087] = -13'h000f;
         mem[2088] =  13'h007f;
         mem[2089] =  13'h0067;
         mem[2090] = -13'h0073;
         mem[2091] =  13'h0095;
         mem[2092] = -13'h0128;
         mem[2093] = -13'h00aa;
         mem[2094] =  13'h00c3;
         mem[2095] =  13'h010d;
         mem[2096] =  13'h0038;
         mem[2097] = -13'h0071;
         mem[2098] = -13'h0041;
         mem[2099] =  13'h012f;
         mem[2100] = -13'h0003;
         mem[2101] =  13'h0049;
         mem[2102] = -13'h000a;
         mem[2103] = -13'h0025;
         mem[2104] =  13'h00c9;
         mem[2105] = -13'h007d;
         mem[2106] =  13'h019a;
         mem[2107] =  13'h000d;
         mem[2108] =  13'h0091;
         mem[2109] =  13'h0001;
         mem[2110] =  13'h0067;
         mem[2111] = -13'h0015;
         mem[2112] =  13'h0006;
         mem[2113] = -13'h0042;
         mem[2114] = -13'h0079;
         mem[2115] = -13'h0006;
         mem[2116] = -13'h00dd;
         mem[2117] = -13'h010f;
         mem[2118] =  13'h0072;
         mem[2119] =  13'h0076;
         mem[2120] = -13'h0053;
         mem[2121] =  13'h0032;
         mem[2122] =  13'h00b1;
         mem[2123] =  13'h02fa;
         mem[2124] =  13'h0082;
         mem[2125] =  13'h0039;
         mem[2126] = -13'h0019;
         mem[2127] = -13'h0016;
         mem[2128] =  13'h0044;
         mem[2129] =  13'h006a;
         mem[2130] = -13'h006d;
         mem[2131] = -13'h0045;
         mem[2132] =  13'h0018;
         mem[2133] = -13'h000b;
         mem[2134] = -13'h00b3;
         mem[2135] =  13'h00d3;
         mem[2136] =  13'h0021;
         mem[2137] = -13'h00d8;
         mem[2138] =  13'h00d7;
         mem[2139] = -13'h0033;
         mem[2140] =  13'h002f;
         mem[2141] = -13'h0061;
         mem[2142] = -13'h00fc;
         mem[2143] = -13'h0007;
         mem[2144] =  13'h0090;
         mem[2145] = -13'h004b;
         mem[2146] = -13'h009d;
         mem[2147] =  13'h0198;
         mem[2148] =  13'h0159;
         mem[2149] =  13'h00a4;
         mem[2150] =  13'h00f1;
         mem[2151] =  13'h0264;
         mem[2152] =  13'h0002;
         mem[2153] = -13'h0088;
         mem[2154] =  13'h0026;
         mem[2155] =  13'h00b0;
         mem[2156] = -13'h0114;
         mem[2157] = -13'h04fc;
         mem[2158] =  13'h0079;
         mem[2159] =  13'h002b;
         mem[2160] = -13'h0076;
         mem[2161] = -13'h0017;
         mem[2162] =  13'h0074;
         mem[2163] = -13'h0076;
         mem[2164] =  13'h0066;
         mem[2165] =  13'h0031;
         mem[2166] = -13'h00ae;
         mem[2167] =  13'h002a;
         mem[2168] = -13'h011b;
         mem[2169] = -13'h0013;
         mem[2170] = -13'h0039;
         mem[2171] = -13'h003e;
         mem[2172] = -13'h0029;
         mem[2173] = -13'h00d0;
         mem[2174] =  13'h007d;
         mem[2175] = -13'h002d;
         mem[2176] = -13'h0019;
         mem[2177] =  13'h0141;
         mem[2178] = -13'h0029;
         mem[2179] =  13'h007f;
         mem[2180] =  13'h00a4;
         mem[2181] =  13'h0042;
         mem[2182] = -13'h00ba;
         mem[2183] = -13'h004a;
         mem[2184] = -13'h0039;
         mem[2185] = -13'h009e;
         mem[2186] =  13'h0081;
         mem[2187] = -13'h002c;
         mem[2188] =  13'h0031;
         mem[2189] =  13'h0121;
         mem[2190] =  13'h0880;
         mem[2191] = -13'h003c;
         mem[2192] = -13'h0009;
         mem[2193] =  13'h00cc;
         mem[2194] = -13'h00c3;
         mem[2195] = -13'h0176;
         mem[2196] =  13'h009b;
         mem[2197] = -13'h003f;
         mem[2198] = -13'h003f;
         mem[2199] = -13'h00eb;
         mem[2200] = -13'h0018;
         mem[2201] = -13'h011e;
         mem[2202] = -13'h0066;
         mem[2203] =  13'h0046;
         mem[2204] = -13'h00b5;
         mem[2205] =  13'h00b4;
         mem[2206] =  13'h0041;
         mem[2207] = -13'h017b;
         mem[2208] =  13'h0122;
         mem[2209] =  13'h00ec;
         mem[2210] = -13'h0043;
         mem[2211] =  13'h0062;
         mem[2212] =  13'h0033;
         mem[2213] = -13'h00de;
         mem[2214] = -13'h0036;
         mem[2215] =  13'h0019;
         mem[2216] =  13'h0076;
         mem[2217] = -13'h005a;
         mem[2218] =  13'h0015;
         mem[2219] =  13'h0160;
         mem[2220] = -13'h0023;
         mem[2221] =  13'h001b;
         mem[2222] = -13'h001a;
         mem[2223] =  13'h0024;
         mem[2224] =  13'h000d;
         mem[2225] =  13'h00a9;
         mem[2226] = -13'h001b;
         mem[2227] =  13'h007d;
         mem[2228] = -13'h001e;
         mem[2229] =  13'h016c;
         mem[2230] =  13'h001d;
         mem[2231] = -13'h004a;
         mem[2232] = -13'h0069;
         mem[2233] =  13'h01bf;
         mem[2234] = -13'h002e;
         mem[2235] = -13'h00eb;
         mem[2236] =  13'h01a4;
         mem[2237] =  13'h006e;
         mem[2238] = -13'h0037;
         mem[2239] = -13'h0525;
         mem[2240] =  13'h0345;
         mem[2241] = -13'h0120;
         mem[2242] =  13'h009a;
         mem[2243] = -13'h011f;
         mem[2244] =  13'h0102;
         mem[2245] =  13'h0095;
         mem[2246] =  13'h0010;
         mem[2247] = -13'h00c9;
         mem[2248] = -13'h0125;
         mem[2249] = -13'h009b;
         mem[2250] = -13'h000c;
         mem[2251] =  13'h004f;
         mem[2252] =  13'h002e;
         mem[2253] = -13'h0089;
         mem[2254] =  13'h0178;
         mem[2255] =  13'h000f;
         mem[2256] =  13'h0034;
         mem[2257] = -13'h024a;
         mem[2258] = -13'h018c;
         mem[2259] = -13'h0024;
         mem[2260] =  13'h0041;
         mem[2261] =  13'h0120;
         mem[2262] = -13'h009b;
         mem[2263] =  13'h0841;
         mem[2264] = -13'h0086;
         mem[2265] = -13'h0094;
         mem[2266] =  13'h001b;
         mem[2267] = -13'h0042;
         mem[2268] =  13'h0022;
         mem[2269] = -13'h0233;
         mem[2270] =  13'h02d4;
         mem[2271] =  13'h0020;
         mem[2272] =  13'h01c1;
         mem[2273] = -13'h007c;
         mem[2274] = -13'h005e;
         mem[2275] = -13'h000c;
         mem[2276] = -13'h0088;
         mem[2277] =  13'h0036;
         mem[2278] =  13'h003c;
         mem[2279] = -13'h0036;
         mem[2280] = -13'h0042;
         mem[2281] = -13'h0076;
         mem[2282] = -13'h019f;
         mem[2283] =  13'h009a;
         mem[2284] = -13'h0491;
         mem[2285] =  13'h0275;
         mem[2286] =  13'h0000;
         mem[2287] = -13'h0054;
         mem[2288] =  13'h0099;
         mem[2289] =  13'h00ea;
         mem[2290] =  13'h0014;
         mem[2291] = -13'h00df;
         mem[2292] =  13'h0067;
         mem[2293] =  13'h0063;
         mem[2294] =  13'h0093;
         mem[2295] = -13'h0199;
         mem[2296] =  13'h0159;
         mem[2297] =  13'h0041;
         mem[2298] =  13'h008a;
         mem[2299] = -13'h00fd;
         mem[2300] =  13'h011e;
         mem[2301] = -13'h0072;
         mem[2302] = -13'h0034;
         mem[2303] =  13'h0058;
         mem[2304] =  13'h019b;
         mem[2305] =  13'h006a;
         mem[2306] =  13'h0074;
         mem[2307] =  13'h009e;
         mem[2308] = -13'h00be;
         mem[2309] = -13'h00af;
         mem[2310] =  13'h000f;
         mem[2311] =  13'h00ad;
         mem[2312] =  13'h0050;
         mem[2313] =  13'h0003;
         mem[2314] = -13'h0011;
         mem[2315] =  13'h0045;
         mem[2316] =  13'h0093;
         mem[2317] = -13'h0122;
         mem[2318] = -13'h0102;
         mem[2319] =  13'h0079;
         mem[2320] =  13'h009b;
         mem[2321] = -13'h0088;
         mem[2322] = -13'h0081;
         mem[2323] =  13'h0004;
         mem[2324] = -13'h0125;
         mem[2325] = -13'h014c;
         mem[2326] =  13'h0012;
         mem[2327] = -13'h00ac;
         mem[2328] = -13'h010c;
         mem[2329] =  13'h004a;
         mem[2330] = -13'h00d3;
         mem[2331] = -13'h00c1;
         mem[2332] =  13'h0047;
         mem[2333] = -13'h0067;
         mem[2334] = -13'h00a6;
         mem[2335] = -13'h009a;
         mem[2336] = -13'h0036;
         mem[2337] =  13'h0000;
         mem[2338] = -13'h002e;
         mem[2339] =  13'h0098;
         mem[2340] =  13'h000d;
         mem[2341] = -13'h005c;
         mem[2342] =  13'h005f;
         mem[2343] = -13'h0039;
         mem[2344] =  13'h001e;
         mem[2345] = -13'h002f;
         mem[2346] =  13'h00d7;
         mem[2347] =  13'h00d7;
         mem[2348] = -13'h0030;
         mem[2349] =  13'h0188;
         mem[2350] = -13'h0041;
         mem[2351] =  13'h008e;
         mem[2352] =  13'h008e;
         mem[2353] =  13'h0042;
         mem[2354] = -13'h00b5;
         mem[2355] = -13'h0016;
         mem[2356] = -13'h010d;
         mem[2357] = -13'h012c;
         mem[2358] =  13'h0043;
         mem[2359] = -13'h0025;
         mem[2360] =  13'h0018;
         mem[2361] = -13'h0003;
         mem[2362] =  13'h0349;
         mem[2363] = -13'h0045;
         mem[2364] = -13'h004e;
         mem[2365] = -13'h006a;
         mem[2366] = -13'h0059;
         mem[2367] = -13'h0062;
         mem[2368] =  13'h00c1;
         mem[2369] = -13'h00bc;
         mem[2370] =  13'h006c;
         mem[2371] = -13'h00c7;
         mem[2372] = -13'h004c;
         mem[2373] =  13'h0033;
         mem[2374] = -13'h0004;
         mem[2375] = -13'h00c9;
         mem[2376] = -13'h0047;
         mem[2377] = -13'h003c;
         mem[2378] = -13'h03aa;
         mem[2379] = -13'h0208;
         mem[2380] =  13'h002a;
         mem[2381] =  13'h001c;
         mem[2382] =  13'h04a4;
         mem[2383] = -13'h03cf;
         mem[2384] =  13'h00ff;
         mem[2385] =  13'h0013;
         mem[2386] = -13'h0071;
         mem[2387] = -13'h0045;
         mem[2388] = -13'h00cb;
         mem[2389] = -13'h0132;
         mem[2390] =  13'h0083;
         mem[2391] = -13'h0182;
         mem[2392] = -13'h003f;
         mem[2393] = -13'h0010;
         mem[2394] =  13'h000c;
         mem[2395] = -13'h0029;
         mem[2396] = -13'h009e;
         mem[2397] =  13'h008d;
         mem[2398] = -13'h0013;
         mem[2399] =  13'h0002;
         mem[2400] =  13'h0090;
         mem[2401] = -13'h0060;
         mem[2402] = -13'h0007;
         mem[2403] = -13'h0044;
         mem[2404] =  13'h0a91;
         mem[2405] =  13'h01c1;
         mem[2406] =  13'h0037;
         mem[2407] = -13'h005d;
         mem[2408] = -13'h014f;
         mem[2409] = -13'h00d7;
         mem[2410] = -13'h0067;
         mem[2411] = -13'h00b3;
         mem[2412] = -13'h004a;
         mem[2413] =  13'h0060;
         mem[2414] =  13'h008c;
         mem[2415] =  13'h0069;
         mem[2416] = -13'h006c;
         mem[2417] =  13'h00f9;
         mem[2418] =  13'h0250;
         mem[2419] =  13'h00da;
         mem[2420] =  13'h002e;
         mem[2421] = -13'h0009;
         mem[2422] = -13'h0079;
         mem[2423] =  13'h006f;
         mem[2424] = -13'h000e;
         mem[2425] = -13'h0033;
         mem[2426] = -13'h016b;
         mem[2427] = -13'h004e;
         mem[2428] = -13'h0044;
         mem[2429] =  13'h0034;
         mem[2430] = -13'h0037;
         mem[2431] =  13'h004d;
         mem[2432] = -13'h001a;
         mem[2433] = -13'h0063;
         mem[2434] = -13'h0079;
         mem[2435] =  13'h0014;
         mem[2436] = -13'h0017;
         mem[2437] =  13'h0044;
         mem[2438] =  13'h009c;
         mem[2439] = -13'h00e9;
         mem[2440] = -13'h00dc;
         mem[2441] = -13'h000a;
         mem[2442] =  13'h04c1;
         mem[2443] = -13'h016c;
         mem[2444] = -13'h00e6;
         mem[2445] =  13'h0097;
         mem[2446] = -13'h0022;
         mem[2447] = -13'h0009;
         mem[2448] = -13'h0125;
         mem[2449] =  13'h0015;
         mem[2450] = -13'h0019;
         mem[2451] =  13'h003f;
         mem[2452] =  13'h006a;
         mem[2453] = -13'h0031;
         mem[2454] = -13'h0115;
         mem[2455] = -13'h003c;
         mem[2456] =  13'h0066;
         mem[2457] =  13'h004d;
         mem[2458] = -13'h0057;
         mem[2459] =  13'h0026;
         mem[2460] =  13'h03ac;
         mem[2461] = -13'h009b;
         mem[2462] = -13'h0037;
         mem[2463] =  13'h0094;
         mem[2464] =  13'h001b;
         mem[2465] =  13'h018b;
         mem[2466] = -13'h0092;
         mem[2467] =  13'h002c;
         mem[2468] =  13'h0144;
         mem[2469] =  13'h0086;
         mem[2470] = -13'h0071;
         mem[2471] = -13'h0010;
         mem[2472] =  13'h001e;
         mem[2473] =  13'h01cb;
         mem[2474] = -13'h01e6;
         mem[2475] = -13'h00aa;
         mem[2476] = -13'h0072;
         mem[2477] = -13'h0200;
         mem[2478] =  13'h03c9;
         mem[2479] = -13'h0078;
         mem[2480] =  13'h009a;
         mem[2481] =  13'h0127;
         mem[2482] =  13'h0028;
         mem[2483] =  13'h00d5;
         mem[2484] = -13'h00b3;
         mem[2485] = -13'h009d;
         mem[2486] = -13'h0194;
         mem[2487] = -13'h01f3;
         mem[2488] = -13'h01ea;
         mem[2489] =  13'h007e;
         mem[2490] =  13'h002c;
         mem[2491] =  13'h00e8;
         mem[2492] =  13'h0004;
         mem[2493] = -13'h0073;
         mem[2494] = -13'h028f;
         mem[2495] =  13'h0014;
         mem[2496] =  13'h00c0;
         mem[2497] =  13'h0063;
         mem[2498] =  13'h011f;
         mem[2499] =  13'h0028;
         mem[2500] = -13'h00e6;
         mem[2501] =  13'h01c1;
         mem[2502] =  13'h0055;
         mem[2503] =  13'h008f;
         mem[2504] =  13'h00a3;
         mem[2505] = -13'h0013;
         mem[2506] =  13'h0009;
         mem[2507] =  13'h0067;
         mem[2508] = -13'h0083;
         mem[2509] =  13'h0134;
         mem[2510] = -13'h004b;
         mem[2511] = -13'h0034;
         mem[2512] = -13'h006c;
         mem[2513] =  13'h005a;
         mem[2514] =  13'h0258;
         mem[2515] =  13'h000e;
         mem[2516] =  13'h0026;
         mem[2517] = -13'h0023;
         mem[2518] = -13'h00a0;
         mem[2519] =  13'h0065;
         mem[2520] = -13'h008f;
         mem[2521] = -13'h004b;
         mem[2522] = -13'h0037;
         mem[2523] =  13'h0019;
         mem[2524] = -13'h004b;
         mem[2525] =  13'h003a;
         mem[2526] = -13'h0085;
         mem[2527] = -13'h000a;
         mem[2528] = -13'h0003;
         mem[2529] =  13'h00c2;
         mem[2530] = -13'h001c;
         mem[2531] = -13'h00b0;
         mem[2532] =  13'h0054;
         mem[2533] = -13'h005b;
         mem[2534] =  13'h00cc;
         mem[2535] =  13'h00fd;
         mem[2536] = -13'h00ab;
         mem[2537] = -13'h000d;
         mem[2538] =  13'h0063;
         mem[2539] = -13'h0046;
         mem[2540] = -13'h0010;
         mem[2541] = -13'h003a;
         mem[2542] = -13'h0025;
         mem[2543] = -13'h01fa;
         mem[2544] = -13'h0150;
         mem[2545] =  13'h010c;
         mem[2546] = -13'h0081;
         mem[2547] = -13'h0146;
         mem[2548] = -13'h004d;
         mem[2549] = -13'h0014;
         mem[2550] = -13'h0032;
         mem[2551] =  13'h0005;
         mem[2552] =  13'h0079;
         mem[2553] =  13'h0073;
         mem[2554] =  13'h007c;
         mem[2555] = -13'h0046;
         mem[2556] = -13'h0158;
         mem[2557] =  13'h001e;
         mem[2558] =  13'h00e7;
         mem[2559] = -13'h0015;
         mem[2560] = -13'h003d;
         mem[2561] =  13'h00e0;
         mem[2562] = -13'h0050;
         mem[2563] = -13'h0113;
         mem[2564] = -13'h003a;
         mem[2565] =  13'h007a;
         mem[2566] =  13'h00d4;
         mem[2567] =  13'h00a8;
         mem[2568] = -13'h020e;
         mem[2569] =  13'h0009;
         mem[2570] =  13'h001f;
         mem[2571] =  13'h00ba;
         mem[2572] = -13'h0142;
         mem[2573] =  13'h0020;
         mem[2574] = -13'h0037;
         mem[2575] =  13'h0076;
         mem[2576] = -13'h0070;
         mem[2577] = -13'h012a;
         mem[2578] = -13'h0039;
         mem[2579] =  13'h00b1;
         mem[2580] =  13'h0078;
         mem[2581] = -13'h0082;
         mem[2582] =  13'h009b;
         mem[2583] = -13'h005b;
         mem[2584] =  13'h00f1;
         mem[2585] =  13'h007f;
         mem[2586] =  13'h0099;
         mem[2587] = -13'h0055;
         mem[2588] = -13'h0068;
         mem[2589] = -13'h001d;
         mem[2590] = -13'h00d0;
         mem[2591] = -13'h0054;
         mem[2592] =  13'h002b;
         mem[2593] =  13'h0082;
         mem[2594] = -13'h0061;
         mem[2595] = -13'h0018;
         mem[2596] =  13'h0061;
         mem[2597] =  13'h0072;
         mem[2598] =  13'h003b;
         mem[2599] =  13'h01bd;
         mem[2600] = -13'h0039;
         mem[2601] =  13'h0010;
         mem[2602] = -13'h0014;
         mem[2603] = -13'h015c;
         mem[2604] =  13'h0008;
         mem[2605] =  13'h05d2;
         mem[2606] =  13'h0388;
         mem[2607] = -13'h0042;
         mem[2608] = -13'h00c5;
         mem[2609] =  13'h0047;
         mem[2610] = -13'h008c;
         mem[2611] = -13'h0012;
         mem[2612] =  13'h0210;
         mem[2613] =  13'h007c;
         mem[2614] =  13'h00b4;
         mem[2615] =  13'h000c;
         mem[2616] = -13'h006b;
         mem[2617] = -13'h0072;
         mem[2618] =  13'h0030;
         mem[2619] =  13'h0006;
         mem[2620] = -13'h000e;
         mem[2621] = -13'h0081;
         mem[2622] = -13'h0083;
         mem[2623] =  13'h027c;
         mem[2624] =  13'h0168;
         mem[2625] = -13'h0006;
         mem[2626] =  13'h0026;
         mem[2627] =  13'h0098;
         mem[2628] =  13'h0148;
         mem[2629] = -13'h0003;
         mem[2630] = -13'h0014;
         mem[2631] =  13'h01e9;
         mem[2632] = -13'h0012;
         mem[2633] = -13'h0079;
         mem[2634] =  13'h006d;
         mem[2635] =  13'h00b5;
         mem[2636] = -13'h0063;
         mem[2637] =  13'h0050;
         mem[2638] =  13'h0016;
         mem[2639] = -13'h03b6;
         mem[2640] = -13'h0068;
         mem[2641] = -13'h001a;
         mem[2642] =  13'h0010;
         mem[2643] = -13'h0092;
         mem[2644] = -13'h003a;
         mem[2645] = -13'h0205;
         mem[2646] =  13'h0119;
         mem[2647] =  13'h015f;
         mem[2648] =  13'h003f;
         mem[2649] =  13'h014c;
         mem[2650] =  13'h004b;
         mem[2651] = -13'h0161;
         mem[2652] =  13'h0128;
         mem[2653] = -13'h0140;
         mem[2654] =  13'h018c;
         mem[2655] = -13'h00a3;
         mem[2656] = -13'h0027;
         mem[2657] =  13'h0001;
         mem[2658] =  13'h0031;
         mem[2659] = -13'h0055;
         mem[2660] =  13'h00ed;
         mem[2661] =  13'h0000;
         mem[2662] = -13'h0046;
         mem[2663] =  13'h007d;
         mem[2664] = -13'h0003;
         mem[2665] =  13'h0168;
         mem[2666] = -13'h009f;
         mem[2667] =  13'h0148;
         mem[2668] =  13'h00a1;
         mem[2669] =  13'h0054;
         mem[2670] = -13'h0112;
         mem[2671] =  13'h00bf;
         mem[2672] =  13'h0141;
         mem[2673] =  13'h010f;
         mem[2674] =  13'h007b;
         mem[2675] =  13'h0046;
         mem[2676] =  13'h0052;
         mem[2677] =  13'h0087;
         mem[2678] = -13'h003c;
         mem[2679] = -13'h002a;
         mem[2680] = -13'h0075;
         mem[2681] = -13'h0013;
         mem[2682] =  13'h0526;
         mem[2683] = -13'h0045;
         mem[2684] = -13'h001e;
         mem[2685] = -13'h007a;
         mem[2686] = -13'h002e;
         mem[2687] =  13'h0013;
         mem[2688] =  13'h0014;
         mem[2689] =  13'h0318;
         mem[2690] =  13'h0016;
         mem[2691] = -13'h0117;
         mem[2692] = -13'h008f;
         mem[2693] =  13'h0014;
         mem[2694] =  13'h0186;
         mem[2695] = -13'h0101;
         mem[2696] = -13'h02b9;
         mem[2697] =  13'h002b;
         mem[2698] = -13'h00aa;
         mem[2699] =  13'h0208;
         mem[2700] =  13'h0152;
         mem[2701] =  13'h015d;
         mem[2702] =  13'h00e3;
         mem[2703] =  13'h0012;
         mem[2704] =  13'h0035;
         mem[2705] =  13'h00ed;
         mem[2706] = -13'h005d;
         mem[2707] =  13'h00c5;
         mem[2708] =  13'h0069;
         mem[2709] =  13'h001c;
         mem[2710] = -13'h008d;
         mem[2711] =  13'h0078;
         mem[2712] = -13'h0009;
         mem[2713] = -13'h0188;
         mem[2714] =  13'h0044;
         mem[2715] =  13'h006a;
         mem[2716] =  13'h0001;
         mem[2717] = -13'h001b;
         mem[2718] =  13'h004d;
         mem[2719] =  13'h0000;
         mem[2720] = -13'h0138;
         mem[2721] =  13'h00cd;
         mem[2722] = -13'h000b;
         mem[2723] =  13'h0042;
         mem[2724] =  13'h009a;
         mem[2725] = -13'h0032;
         mem[2726] =  13'h00ed;
         mem[2727] =  13'h0013;
         mem[2728] =  13'h00bb;
         mem[2729] =  13'h0057;
         mem[2730] =  13'h0282;
         mem[2731] = -13'h002a;
         mem[2732] =  13'h0009;
         mem[2733] = -13'h005f;
         mem[2734] = -13'h001c;
         mem[2735] = -13'h008c;
         mem[2736] = -13'h0056;
         mem[2737] =  13'h0008;
         mem[2738] = -13'h0011;
         mem[2739] = -13'h003a;
         mem[2740] = -13'h0021;
         mem[2741] = -13'h0026;
         mem[2742] = -13'h009b;
         mem[2743] =  13'h0013;
         mem[2744] = -13'h0012;
         mem[2745] =  13'h0015;
         mem[2746] = -13'h0027;
         mem[2747] =  13'h00b8;
         mem[2748] =  13'h003a;
         mem[2749] =  13'h029e;
         mem[2750] =  13'h000a;
         mem[2751] = -13'h000f;
         mem[2752] = -13'h0067;
         mem[2753] = -13'h004f;
         mem[2754] =  13'h003b;
         mem[2755] =  13'h00d3;
         mem[2756] = -13'h009b;
         mem[2757] = -13'h0079;
         mem[2758] = -13'h00a0;
         mem[2759] = -13'h0077;
         mem[2760] = -13'h0156;
         mem[2761] =  13'h06b8;
         mem[2762] =  13'h00f5;
         mem[2763] = -13'h004d;
         mem[2764] = -13'h0018;
         mem[2765] = -13'h00ee;
         mem[2766] = -13'h0032;
         mem[2767] =  13'h00be;
         mem[2768] =  13'h0004;
         mem[2769] = -13'h016b;
         mem[2770] = -13'h005e;
         mem[2771] =  13'h00b0;
         mem[2772] =  13'h0000;
         mem[2773] =  13'h0024;
         mem[2774] = -13'h0048;
         mem[2775] =  13'h0019;
         mem[2776] =  13'h005d;
         mem[2777] = -13'h0058;
         mem[2778] =  13'h00fc;
         mem[2779] = -13'h013f;
         mem[2780] =  13'h002e;
         mem[2781] = -13'h0068;
         mem[2782] = -13'h009b;
         mem[2783] =  13'h0028;
         mem[2784] = -13'h0038;
         mem[2785] =  13'h0022;
         mem[2786] = -13'h0124;
         mem[2787] =  13'h0028;
         mem[2788] =  13'h01c2;
         mem[2789] =  13'h0090;
         mem[2790] = -13'h01c9;
         mem[2791] = -13'h01d1;
         mem[2792] =  13'h0044;
         mem[2793] = -13'h0020;
         mem[2794] = -13'h0087;
         mem[2795] =  13'h0033;
         mem[2796] = -13'h00ac;
         mem[2797] =  13'h0067;
         mem[2798] = -13'h0063;
         mem[2799] = -13'h0032;
         mem[2800] = -13'h01d2;
         mem[2801] = -13'h015b;
         mem[2802] = -13'h0064;
         mem[2803] = -13'h0024;
         mem[2804] =  13'h002d;
         mem[2805] = -13'h0078;
         mem[2806] =  13'h001a;
         mem[2807] =  13'h0039;
         mem[2808] = -13'h0036;
         mem[2809] =  13'h048c;
         mem[2810] = -13'h03cb;
         mem[2811] = -13'h01c9;
         mem[2812] =  13'h020b;
         mem[2813] = -13'h0101;
         mem[2814] =  13'h0047;
         mem[2815] =  13'h0005;
         mem[2816] =  13'h0070;
         mem[2817] = -13'h00b2;
         mem[2818] =  13'h002d;
         mem[2819] =  13'h0055;
         mem[2820] = -13'h005b;
         mem[2821] =  13'h0085;
         mem[2822] =  13'h0032;
         mem[2823] =  13'h0022;
         mem[2824] =  13'h0099;
         mem[2825] = -13'h0039;
         mem[2826] =  13'h00e9;
         mem[2827] =  13'h0014;
         mem[2828] = -13'h0064;
         mem[2829] = -13'h002e;
         mem[2830] =  13'h008d;
         mem[2831] =  13'h0063;
         mem[2832] = -13'h0020;
         mem[2833] =  13'h008f;
         mem[2834] =  13'h0012;
         mem[2835] = -13'h0154;
         mem[2836] = -13'h0039;
         mem[2837] =  13'h0005;
         mem[2838] = -13'h0044;
         mem[2839] = -13'h013a;
         mem[2840] = -13'h03c9;
         mem[2841] = -13'h019b;
         mem[2842] =  13'h0005;
         mem[2843] =  13'h005a;
         mem[2844] = -13'h01cc;
         mem[2845] =  13'h0043;
         mem[2846] =  13'h0116;
         mem[2847] =  13'h0041;
         mem[2848] =  13'h0013;
         mem[2849] =  13'h001b;
         mem[2850] =  13'h0013;
         mem[2851] =  13'h000a;
         mem[2852] =  13'h000b;
         mem[2853] = -13'h007b;
         mem[2854] =  13'h003a;
         mem[2855] = -13'h00f7;
         mem[2856] = -13'h0051;
         mem[2857] =  13'h007f;
         mem[2858] =  13'h004a;
         mem[2859] =  13'h0004;
         mem[2860] = -13'h0096;
         mem[2861] =  13'h0031;
         mem[2862] =  13'h0132;
         mem[2863] = -13'h03c1;
         mem[2864] =  13'h0241;
         mem[2865] =  13'h0019;
         mem[2866] = -13'h00ea;
         mem[2867] = -13'h00e2;
         mem[2868] = -13'h0058;
         mem[2869] =  13'h0069;
         mem[2870] = -13'h0035;
         mem[2871] =  13'h0009;
         mem[2872] =  13'h0024;
         mem[2873] = -13'h0024;
         mem[2874] =  13'h0010;
         mem[2875] =  13'h0066;
         mem[2876] = -13'h0018;
         mem[2877] =  13'h0011;
         mem[2878] = -13'h008a;
         mem[2879] =  13'h00b6;
         mem[2880] = -13'h00a7;
         mem[2881] =  13'h00a1;
         mem[2882] = -13'h0120;
         mem[2883] =  13'h0092;
         mem[2884] = -13'h00af;
         mem[2885] = -13'h0056;
         mem[2886] = -13'h0284;
         mem[2887] =  13'h0020;
         mem[2888] =  13'h0060;
         mem[2889] =  13'h0131;
         mem[2890] = -13'h0002;
         mem[2891] = -13'h0042;
         mem[2892] = -13'h0087;
         mem[2893] =  13'h00c7;
         mem[2894] =  13'h0009;
         mem[2895] =  13'h00b9;
         mem[2896] =  13'h01b6;
         mem[2897] = -13'h00a5;
         mem[2898] =  13'h0082;
         mem[2899] = -13'h00eb;
         mem[2900] =  13'h0037;
         mem[2901] =  13'h0124;
         mem[2902] = -13'h003d;
         mem[2903] = -13'h0029;
         mem[2904] =  13'h000f;
         mem[2905] =  13'h0042;
         mem[2906] = -13'h00a4;
         mem[2907] =  13'h006e;
         mem[2908] =  13'h00d6;
         mem[2909] = -13'h004e;
         mem[2910] = -13'h000f;
         mem[2911] =  13'h0136;
         mem[2912] = -13'h005a;
     end

endmodule: featureThreshold_rom
