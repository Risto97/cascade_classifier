module passVal_rom
  #(
     parameter W_DATA = 13,
     parameter W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input en1,
     input [W_ADDR-1:0] addr1,
     output reg [W_DATA-1:0] data1

     );

     (* rom_style = "block" *)

     always_ff @(posedge clk)
        begin
           if(en1)
             case(addr1)
               12'b000000000000: data1 <= -13'h0237;
               12'b000000000001: data1 <= 13'h0153;
               12'b000000000010: data1 <= 13'h0110;
               12'b000000000011: data1 <= 13'h012d;
               12'b000000000100: data1 <= 13'h0142;
               12'b000000000101: data1 <= -13'h01df;
               12'b000000000110: data1 <= 13'h0070;
               12'b000000000111: data1 <= 13'h0071;
               12'b000000001000: data1 <= 13'h00da;
               12'b000000001001: data1 <= -13'h0192;
               12'b000000001010: data1 <= 13'h012e;
               12'b000000001011: data1 <= 13'h00b3;
               12'b000000001100: data1 <= 13'h01ba;
               12'b000000001101: data1 <= -13'h022e;
               12'b000000001110: data1 <= 13'h0074;
               12'b000000001111: data1 <= 13'h0089;
               12'b000000010000: data1 <= 13'h00ee;
               12'b000000010001: data1 <= -13'h00a9;
               12'b000000010010: data1 <= -13'h004c;
               12'b000000010011: data1 <= 13'h015b;
               12'b000000010100: data1 <= -13'h0032;
               12'b000000010101: data1 <= -13'h0087;
               12'b000000010110: data1 <= 13'h0124;
               12'b000000010111: data1 <= 13'h00c5;
               12'b000000011000: data1 <= -13'h0183;
               12'b000000011001: data1 <= 13'h0177;
               12'b000000011010: data1 <= 13'h0100;
               12'b000000011011: data1 <= -13'h0198;
               12'b000000011100: data1 <= 13'h00d4;
               12'b000000011101: data1 <= 13'h006c;
               12'b000000011110: data1 <= 13'h010d;
               12'b000000011111: data1 <= -13'h0158;
               12'b000000100000: data1 <= 13'h0173;
               12'b000000100001: data1 <= 13'h0136;
               12'b000000100010: data1 <= -13'h0075;
               12'b000000100011: data1 <= 13'h0027;
               12'b000000100100: data1 <= -13'h0190;
               12'b000000100101: data1 <= 13'h003b;
               12'b000000100110: data1 <= 13'h0147;
               12'b000000100111: data1 <= -13'h004d;
               12'b000000101000: data1 <= -13'h000d;
               12'b000000101001: data1 <= 13'h0189;
               12'b000000101010: data1 <= 13'h00ef;
               12'b000000101011: data1 <= 13'h00f6;
               12'b000000101100: data1 <= -13'h02f5;
               12'b000000101101: data1 <= -13'h0070;
               12'b000000101110: data1 <= 13'h0066;
               12'b000000101111: data1 <= -13'h02a5;
               12'b000000110000: data1 <= 13'h0048;
               12'b000000110001: data1 <= 13'h003b;
               12'b000000110010: data1 <= 13'h0113;
               12'b000000110011: data1 <= 13'h0019;

endmodule: passVal_rom
