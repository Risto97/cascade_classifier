module rect0_rom
  #(
     W_DATA = 20,
     DEPTH = 2913,
     W_ADDR = 12
     )
    (
     input clk,
     input rst,

     input ena,
     input [W_ADDR-1:0] addra,
     output [W_DATA-1:0] doa
    );

     logic [W_DATA-1:0] mem [DEPTH-1:0];

     always_ff @(posedge clk)
        begin
           if(ena)
              doa = mem[addra];
        end

     initial begin
         mem[0] =  20'h1a989;
         mem[1] =  20'h1a987;
         mem[2] =  20'h39249;
         mem[3] =  20'h72926;
         mem[4] =  20'h20093;
         mem[5] =  20'h20d90;
         mem[6] =  20'h33586;
         mem[7] =  20'h5a48a;
         mem[8] =  20'h010e6;
         mem[9] =  20'h27186;
         mem[10] =  20'h1a987;
         mem[11] =  20'h3266c;
         mem[12] =  20'h0cb03;
         mem[13] =  20'h3a8cf;
         mem[14] =  20'h26dca;
         mem[15] =  20'h015c9;
         mem[16] =  20'h48126;
         mem[17] =  20'h210ca;
         mem[18] =  20'h348ca;
         mem[19] =  20'h1fc89;
         mem[20] =  20'h048cb;
         mem[21] =  20'h25b0d;
         mem[22] =  20'h27cc9;
         mem[23] =  20'h72546;
         mem[24] =  20'h2d1cc;
         mem[25] =  20'h12f03;
         mem[26] =  20'h335e6;
         mem[27] =  20'h27cae;
         mem[28] =  20'h218ca;
         mem[29] =  20'h2706c;
         mem[30] =  20'h84243;
         mem[31] =  20'h26da6;
         mem[32] =  20'h0accf;
         mem[33] =  20'h068cf;
         mem[34] =  20'h3230f;
         mem[35] =  20'h26dcc;
         mem[36] =  20'h4baac;
         mem[37] =  20'h0848a;
         mem[38] =  20'h51e8a;
         mem[39] =  20'h064cd;
         mem[40] =  20'h1188d;
         mem[41] =  20'h1f6d3;
         mem[42] =  20'h1d8c9;
         mem[43] =  20'h12ccb;
         mem[44] =  20'h09489;
         mem[45] =  20'h25a63;
         mem[46] =  20'h09489;
         mem[47] =  20'h08489;
         mem[48] =  20'h209ce;
         mem[49] =  20'h3ee42;
         mem[50] =  20'h5588b;
         mem[51] =  20'h190c9;
         mem[52] =  20'h1a989;
         mem[53] =  20'h20d86;
         mem[54] =  20'h06705;
         mem[55] =  20'h3fa46;
         mem[56] =  20'h6ad86;
         mem[57] =  20'h1788d;
         mem[58] =  20'h1308d;
         mem[59] =  20'h06717;
         mem[60] =  20'h2c10c;
         mem[61] =  20'h2f46e;
         mem[62] =  20'h4be06;
         mem[63] =  20'h27186;
         mem[64] =  20'h2dccc;
         mem[65] =  20'h61926;
         mem[66] =  20'h6aa43;
         mem[67] =  20'h1a20c;
         mem[68] =  20'h06494;
         mem[69] =  20'h00e42;
         mem[70] =  20'h1fa8e;
         mem[71] =  20'h335cc;
         mem[72] =  20'h584e9;
         mem[73] =  20'h61526;
         mem[74] =  20'h5e126;
         mem[75] =  20'h2850a;
         mem[76] =  20'h209ce;
         mem[77] =  20'h01985;
         mem[78] =  20'h024c9;
         mem[79] =  20'h27cc9;
         mem[80] =  20'h01cc9;
         mem[81] =  20'h280c9;
         mem[82] =  20'h278c9;
         mem[83] =  20'h32e44;
         mem[84] =  20'h01989;
         mem[85] =  20'h00306;
         mem[86] =  20'h2ce0c;
         mem[87] =  20'h284c6;
         mem[88] =  20'h7d303;
         mem[89] =  20'h28489;
         mem[90] =  20'h525e4;
         mem[91] =  20'h28489;
         mem[92] =  20'h27c89;
         mem[93] =  20'h4d4cc;
         mem[94] =  20'h89e42;
         mem[95] =  20'h2e48a;
         mem[96] =  20'h2d50a;
         mem[97] =  20'h27546;
         mem[98] =  20'h57944;
         mem[99] =  20'h72242;
         mem[100] =  20'h06ac3;
         mem[101] =  20'h65a43;
         mem[102] =  20'h198cf;
         mem[103] =  20'h1e08a;
         mem[104] =  20'h1908a;
         mem[105] =  20'h64a86;
         mem[106] =  20'h4b109;
         mem[107] =  20'h030c9;
         mem[108] =  20'h3fcc6;
         mem[109] =  20'h34d86;
         mem[110] =  20'h32186;
         mem[111] =  20'h030c9;
         mem[112] =  20'h018c9;
         mem[113] =  20'h59926;
         mem[114] =  20'h64126;
         mem[115] =  20'h348ca;
         mem[116] =  20'h77983;
         mem[117] =  20'h3f282;
         mem[118] =  20'h38e4c;
         mem[119] =  20'h00e58;
         mem[120] =  20'h26dca;
         mem[121] =  20'h2194c;
         mem[122] =  20'h2058c;
         mem[123] =  20'h58a43;
         mem[124] =  20'h52d08;
         mem[125] =  20'h64e46;
         mem[126] =  20'h000c6;
         mem[127] =  20'h27192;
         mem[128] =  20'h07c8e;
         mem[129] =  20'h0d662;
         mem[130] =  20'h326cd;
         mem[131] =  20'h3a564;
         mem[132] =  20'h4b1ea;
         mem[133] =  20'h67186;
         mem[134] =  20'h64186;
         mem[135] =  20'h0b0ac;
         mem[136] =  20'h0cb04;
         mem[137] =  20'h33984;
         mem[138] =  20'h21126;
         mem[139] =  20'h6c8c6;
         mem[140] =  20'h2becf;
         mem[141] =  20'h07629;
         mem[142] =  20'h210ca;
         mem[143] =  20'h0acc8;
         mem[144] =  20'h064c7;
         mem[145] =  20'h048d6;
         mem[146] =  20'h000d6;
         mem[147] =  20'h2fd10;
         mem[148] =  20'h3f266;
         mem[149] =  20'h3a8cc;
         mem[150] =  20'h5e626;
         mem[151] =  20'h2f46e;
         mem[152] =  20'h26d0a;
         mem[153] =  20'h35d2b;
         mem[154] =  20'h3212b;
         mem[155] =  20'h27952;
         mem[156] =  20'h2d86e;
         mem[157] =  20'h57b08;
         mem[158] =  20'h3ee4e;
         mem[159] =  20'h4e8c6;
         mem[160] =  20'h01d50;
         mem[161] =  20'h02926;
         mem[162] =  20'h13e04;
         mem[163] =  20'h02926;
         mem[164] =  20'h06a84;
         mem[165] =  20'h02926;
         mem[166] =  20'h01526;
         mem[167] =  20'h72946;
         mem[168] =  20'h144c9;
         mem[169] =  20'h14986;
         mem[170] =  20'h3ea43;
         mem[171] =  20'h3eec3;
         mem[172] =  20'h46108;
         mem[173] =  20'h47cc6;
         mem[174] =  20'h464c6;
         mem[175] =  20'h40566;
         mem[176] =  20'h51704;
         mem[177] =  20'h19acc;
         mem[178] =  20'h00a91;
         mem[179] =  20'h03858;
         mem[180] =  20'h02058;
         mem[181] =  20'h09c56;
         mem[182] =  20'h08456;
         mem[183] =  20'h29c72;
         mem[184] =  20'h59126;
         mem[185] =  20'h5ad24;
         mem[186] =  20'h71643;
         mem[187] =  20'h1b512;
         mem[188] =  20'h6a643;
         mem[189] =  20'h0c984;
         mem[190] =  20'h339c6;
         mem[191] =  20'h210c6;
         mem[192] =  20'h21cd0;
         mem[193] =  20'h19530;
         mem[194] =  20'h01649;
         mem[195] =  20'h600a8;
         mem[196] =  20'h05089;
         mem[197] =  20'h00a43;
         mem[198] =  20'h8ae62;
         mem[199] =  20'h00089;
         mem[200] =  20'h26e72;
         mem[201] =  20'h064c9;
         mem[202] =  20'h20dcc;
         mem[203] =  20'h06682;
         mem[204] =  20'h0cec3;
         mem[205] =  20'h328e9;
         mem[206] =  20'h4bac4;
         mem[207] =  20'h4b2c4;
         mem[208] =  20'h2e0cb;
         mem[209] =  20'h08126;
         mem[210] =  20'h0f48a;
         mem[211] =  20'h1a98c;
         mem[212] =  20'h0accf;
         mem[213] =  20'h5ea43;
         mem[214] =  20'h23cc9;
         mem[215] =  20'h1fa06;
         mem[216] =  20'h02cc9;
         mem[217] =  20'h1930e;
         mem[218] =  20'h0348d;
         mem[219] =  20'h01c8d;
         mem[220] =  20'h284c9;
         mem[221] =  20'h2dcc9;
         mem[222] =  20'h6d926;
         mem[223] =  20'h711c6;
         mem[224] =  20'h71644;
         mem[225] =  20'h7d1e4;
         mem[226] =  20'h601e9;
         mem[227] =  20'h1a204;
         mem[228] =  20'h27546;
         mem[229] =  20'h579ea;
         mem[230] =  20'h3a14e;
         mem[231] =  20'h274c9;
         mem[232] =  20'h26643;
         mem[233] =  20'h3ea43;
         mem[234] =  20'h64e44;
         mem[235] =  20'h269c6;
         mem[236] =  20'h03452;
         mem[237] =  20'h02452;
         mem[238] =  20'h2d1ea;
         mem[239] =  20'h7d6a4;
         mem[240] =  20'h21cb2;
         mem[241] =  20'h0cb06;
         mem[242] =  20'h06ac8;
         mem[243] =  20'h011e9;
         mem[244] =  20'h00313;
         mem[245] =  20'h83e43;
         mem[246] =  20'h2e144;
         mem[247] =  20'h2d144;
         mem[248] =  20'h364d0;
         mem[249] =  20'h5e284;
         mem[250] =  20'h61546;
         mem[251] =  20'h00e09;
         mem[252] =  20'h294ef;
         mem[253] =  20'h088cd;
         mem[254] =  20'h10cce;
         mem[255] =  20'h5858a;
         mem[256] =  20'h27546;
         mem[257] =  20'h0ccce;
         mem[258] =  20'h1b8ac;
         mem[259] =  20'h6a705;
         mem[260] =  20'h2f8ac;
         mem[261] =  20'h070cc;
         mem[262] =  20'h544c6;
         mem[263] =  20'h52cc6;
         mem[264] =  20'h29070;
         mem[265] =  20'h4b5a6;
         mem[266] =  20'h09889;
         mem[267] =  20'h01d26;
         mem[268] =  20'h0f8c9;
         mem[269] =  20'h0e0c9;
         mem[270] =  20'h72186;
         mem[271] =  20'h274c9;
         mem[272] =  20'h2d983;
         mem[273] =  20'h14d15;
         mem[274] =  20'h1ad4c;
         mem[275] =  20'h064c9;
         mem[276] =  20'h10454;
         mem[277] =  20'h12cc9;
         mem[278] =  20'h16855;
         mem[279] =  20'h01c57;
         mem[280] =  20'h35d24;
         mem[281] =  20'h32124;
         mem[282] =  20'h59926;
         mem[283] =  20'h57926;
         mem[284] =  20'h3f644;
         mem[285] =  20'h00313;
         mem[286] =  20'h0890c;
         mem[287] =  20'h2808a;
         mem[288] =  20'h3a14c;
         mem[289] =  20'h01473;
         mem[290] =  20'h038ca;
         mem[291] =  20'h008cc;
         mem[292] =  20'h44f02;
         mem[293] =  20'h395a4;
         mem[294] =  20'h344c9;
         mem[295] =  20'h4b204;
         mem[296] =  20'h4f8c9;
         mem[297] =  20'h4b0c9;
         mem[298] =  20'h2dd44;
         mem[299] =  20'h2dcc9;
         mem[300] =  20'h02cc9;
         mem[301] =  20'h01cc9;
         mem[302] =  20'h15ccf;
         mem[303] =  20'h144cf;
         mem[304] =  20'h10524;
         mem[305] =  20'h3fcc7;
         mem[306] =  20'h59cca;
         mem[307] =  20'h530a8;
         mem[308] =  20'h22c70;
         mem[309] =  20'h6ae43;
         mem[310] =  20'h71e63;
         mem[311] =  20'h024c9;
         mem[312] =  20'h1c072;
         mem[313] =  20'h1b472;
         mem[314] =  20'h13a49;
         mem[315] =  20'h07cce;
         mem[316] =  20'h67126;
         mem[317] =  20'h13290;
         mem[318] =  20'h224cc;
         mem[319] =  20'h0ced0;
         mem[320] =  20'h5a0aa;
         mem[321] =  20'h84243;
         mem[322] =  20'h5a0ca;
         mem[323] =  20'h0cb04;
         mem[324] =  20'h1a989;
         mem[325] =  20'h27185;
         mem[326] =  20'h335cc;
         mem[327] =  20'h5890a;
         mem[328] =  20'h284ae;
         mem[329] =  20'h27470;
         mem[330] =  20'h2ca48;
         mem[331] =  20'h13682;
         mem[332] =  20'h4be66;
         mem[333] =  20'h278c9;
         mem[334] =  20'h298ce;
         mem[335] =  20'h3a0cc;
         mem[336] =  20'h2a0d2;
         mem[337] =  20'h258d2;
         mem[338] =  20'h110c9;
         mem[339] =  20'h715e6;
         mem[340] =  20'h110c9;
         mem[341] =  20'h0c8c9;
         mem[342] =  20'h3fe42;
         mem[343] =  20'h01986;
         mem[344] =  20'h028c9;
         mem[345] =  20'h020c9;
         mem[346] =  20'h4ed26;
         mem[347] =  20'h265a6;
         mem[348] =  20'h4ed26;
         mem[349] =  20'h1fccf;
         mem[350] =  20'h34126;
         mem[351] =  20'h2786e;
         mem[352] =  20'h4ed26;
         mem[353] =  20'h4c144;
         mem[354] =  20'h09893;
         mem[355] =  20'h08093;
         mem[356] =  20'h3ccc9;
         mem[357] =  20'h83a43;
         mem[358] =  20'h54d49;
         mem[359] =  20'h51ac4;
         mem[360] =  20'h26a06;
         mem[361] =  20'h00656;
         mem[362] =  20'h2e50e;
         mem[363] =  20'h190d4;
         mem[364] =  20'h03cc9;
         mem[365] =  20'h00cc9;
         mem[366] =  20'h4eccc;
         mem[367] =  20'h4bccc;
         mem[368] =  20'h4ed26;
         mem[369] =  20'h4b126;
         mem[370] =  20'h58a63;
         mem[371] =  20'h51e63;
         mem[372] =  20'h61546;
         mem[373] =  20'h0194c;
         mem[374] =  20'h0a8cc;
         mem[375] =  20'h068cc;
         mem[376] =  20'h5b8c9;
         mem[377] =  20'h1492c;
         mem[378] =  20'h0948c;
         mem[379] =  20'h011c8;
         mem[380] =  20'h280c9;
         mem[381] =  20'h3f243;
         mem[382] =  20'h61926;
         mem[383] =  20'h066b7;
         mem[384] =  20'h39e24;
         mem[385] =  20'h00572;
         mem[386] =  20'h5f5a6;
         mem[387] =  20'h5dd26;
         mem[388] =  20'h2dde4;
         mem[389] =  20'h4d4c9;
         mem[390] =  20'h33a43;
         mem[391] =  20'h57b04;
         mem[392] =  20'h4286c;
         mem[393] =  20'h12f03;
         mem[394] =  20'h6dd46;
         mem[395] =  20'h51a43;
         mem[396] =  20'h01649;
         mem[397] =  20'h13e09;
         mem[398] =  20'h2346c;
         mem[399] =  20'h2be44;
         mem[400] =  20'h280c9;
         mem[401] =  20'h344ca;
         mem[402] =  20'h600c9;
         mem[403] =  20'h07255;
         mem[404] =  20'h33987;
         mem[405] =  20'h214c9;
         mem[406] =  20'h0cb04;
         mem[407] =  20'h2f4ac;
         mem[408] =  20'h2d0ac;
         mem[409] =  20'h27cc9;
         mem[410] =  20'h064d1;
         mem[411] =  20'h07269;
         mem[412] =  20'h71586;
         mem[413] =  20'h1e093;
         mem[414] =  20'h64147;
         mem[415] =  20'h2dd4c;
         mem[416] =  20'h2d54c;
         mem[417] =  20'h0ed26;
         mem[418] =  20'h7d6a4;
         mem[419] =  20'h4d526;
         mem[420] =  20'h0e526;
         mem[421] =  20'h0348e;
         mem[422] =  20'h01c8e;
         mem[423] =  20'h61526;
         mem[424] =  20'h32a45;
         mem[425] =  20'h174cb;
         mem[426] =  20'h20d6e;
         mem[427] =  20'h1d8c9;
         mem[428] =  20'h27526;
         mem[429] =  20'h1d8c9;
         mem[430] =  20'h190c9;
         mem[431] =  20'h1b524;
         mem[432] =  20'h89a62;
         mem[433] =  20'h5bcc9;
         mem[434] =  20'h57cc9;
         mem[435] =  20'h48489;
         mem[436] =  20'h46489;
         mem[437] =  20'h39247;
         mem[438] =  20'h4d4ca;
         mem[439] =  20'h030c9;
         mem[440] =  20'h018c9;
         mem[441] =  20'h6be43;
         mem[442] =  20'h6aa43;
         mem[443] =  20'h2816c;
         mem[444] =  20'h26dc6;
         mem[445] =  20'h1a5e4;
         mem[446] =  20'h002c2;
         mem[447] =  20'h00318;
         mem[448] =  20'h5e244;
         mem[449] =  20'h33989;
         mem[450] =  20'h4c0ec;
         mem[451] =  20'h0cec6;
         mem[452] =  20'h7e5c3;
         mem[453] =  20'h00310;
         mem[454] =  20'h52244;
         mem[455] =  20'h3f2c2;
         mem[456] =  20'h14568;
         mem[457] =  20'h22cc6;
         mem[458] =  20'h2bf06;
         mem[459] =  20'h0394a;
         mem[460] =  20'h0014a;
         mem[461] =  20'h06704;
         mem[462] =  20'h6a643;
         mem[463] =  20'h5f206;
         mem[464] =  20'h5ea06;
         mem[465] =  20'h65a43;
         mem[466] =  20'h516aa;
         mem[467] =  20'h034d8;
         mem[468] =  20'h1accb;
         mem[469] =  20'h21926;
         mem[470] =  20'h19454;
         mem[471] =  20'h034d8;
         mem[472] =  20'h014d8;
         mem[473] =  20'h2fcce;
         mem[474] =  20'h2cc8c;
         mem[475] =  20'h1f70e;
         mem[476] =  20'h52946;
         mem[477] =  20'h030c9;
         mem[478] =  20'h2c4ce;
         mem[479] =  20'h1052f;
         mem[480] =  20'h0c8c9;
         mem[481] =  20'h0f94e;
         mem[482] =  20'h28452;
         mem[483] =  20'h219e6;
         mem[484] =  20'h278ca;
         mem[485] =  20'h030c9;
         mem[486] =  20'h13927;
         mem[487] =  20'h2d5c3;
         mem[488] =  20'h2d906;
         mem[489] =  20'h2ecec;
         mem[490] =  20'h28092;
         mem[491] =  20'h5b8c9;
         mem[492] =  20'h010cd;
         mem[493] =  20'h0d2a3;
         mem[494] =  20'h1a4ac;
         mem[495] =  20'h1548a;
         mem[496] =  20'h1b0a8;
         mem[497] =  20'h01969;
         mem[498] =  20'h27185;
         mem[499] =  20'h00305;
         mem[500] =  20'h3eee6;
         mem[501] =  20'h84243;
         mem[502] =  20'h266a6;
         mem[503] =  20'h1f4cc;
         mem[504] =  20'h0f08f;
         mem[505] =  20'h2dd0a;
         mem[506] =  20'h2d1ec;
         mem[507] =  20'h6a546;
         mem[508] =  20'h74126;
         mem[509] =  20'h27cd0;
         mem[510] =  20'h74126;
         mem[511] =  20'h70d26;
         mem[512] =  20'h3c126;
         mem[513] =  20'h38526;
         mem[514] =  20'h170c9;
         mem[515] =  20'h6ae43;
         mem[516] =  20'h5eaa6;
         mem[517] =  20'h6c8c6;
         mem[518] =  20'h174c9;
         mem[519] =  20'h12cc9;
         mem[520] =  20'h0120a;
         mem[521] =  20'h00950;
         mem[522] =  20'h03945;
         mem[523] =  20'h00145;
         mem[524] =  20'h174ca;
         mem[525] =  20'h46186;
         mem[526] =  20'h05472;
         mem[527] =  20'h018c9;
         mem[528] =  20'h34127;
         mem[529] =  20'h4cd0a;
         mem[530] =  20'h05472;
         mem[531] =  20'h28089;
         mem[532] =  20'h03d26;
         mem[533] =  20'h0cb03;
         mem[534] =  20'h2e8c9;
         mem[535] =  20'h274ca;
         mem[536] =  20'h094cc;
         mem[537] =  20'h1a98c;
         mem[538] =  20'h16455;
         mem[539] =  20'h07d88;
         mem[540] =  20'h00e48;
         mem[541] =  20'h00e43;
         mem[542] =  20'h51704;
         mem[543] =  20'h21c89;
         mem[544] =  20'h090c9;
         mem[545] =  20'h0e0d6;
         mem[546] =  20'h4290e;
         mem[547] =  20'h19e0f;
         mem[548] =  20'h4290e;
         mem[549] =  20'h3e90e;
         mem[550] =  20'h5a166;
         mem[551] =  20'h2bf09;
         mem[552] =  20'h09890;
         mem[553] =  20'h08090;
         mem[554] =  20'h20a08;
         mem[555] =  20'h384c9;
         mem[556] =  20'h65a43;
         mem[557] =  20'h4bcc9;
         mem[558] =  20'h59926;
         mem[559] =  20'h51d0a;
         mem[560] =  20'h23072;
         mem[561] =  20'h20243;
         mem[562] =  20'h238cb;
         mem[563] =  20'h1f8cb;
         mem[564] =  20'h0b089;
         mem[565] =  20'h06889;
         mem[566] =  20'h5ee49;
         mem[567] =  20'h39d84;
         mem[568] =  20'h10526;
         mem[569] =  20'h0c926;
         mem[570] =  20'h03cd1;
         mem[571] =  20'h00cd1;
         mem[572] =  20'h6c524;
         mem[573] =  20'h20c72;
         mem[574] =  20'h0ddcc;
         mem[575] =  20'h0f06c;
         mem[576] =  20'h2e5cf;
         mem[577] =  20'h2bdcf;
         mem[578] =  20'h03d26;
         mem[579] =  20'h00126;
         mem[580] =  20'h288ce;
         mem[581] =  20'h2e0c9;
         mem[582] =  20'h288cf;
         mem[583] =  20'h270cf;
         mem[584] =  20'h16909;
         mem[585] =  20'h00135;
         mem[586] =  20'h3b10c;
         mem[587] =  20'h2d54c;
         mem[588] =  20'h28092;
         mem[589] =  20'h000c9;
         mem[590] =  20'h58643;
         mem[591] =  20'h5850a;
         mem[592] =  20'h4b304;
         mem[593] =  20'h0c874;
         mem[594] =  20'h67148;
         mem[595] =  20'h64948;
         mem[596] =  20'h01d49;
         mem[597] =  20'h00303;
         mem[598] =  20'h32de4;
         mem[599] =  20'h20d86;
         mem[600] =  20'h529c6;
         mem[601] =  20'h5a48a;
         mem[602] =  20'h258c7;
         mem[603] =  20'h048c6;
         mem[604] =  20'h07243;
         mem[605] =  20'h27dd2;
         mem[606] =  20'h000c6;
         mem[607] =  20'h480c6;
         mem[608] =  20'h7d303;
         mem[609] =  20'h480c7;
         mem[610] =  20'h4c146;
         mem[611] =  20'h480c6;
         mem[612] =  20'h460c7;
         mem[613] =  20'h1ad6c;
         mem[614] =  20'h5f544;
         mem[615] =  20'h038c9;
         mem[616] =  20'h010c9;
         mem[617] =  20'h0f48f;
         mem[618] =  20'h00283;
         mem[619] =  20'h73d46;
         mem[620] =  20'h2c4cb;
         mem[621] =  20'h5a149;
         mem[622] =  20'h0e889;
         mem[623] =  20'h16544;
         mem[624] =  20'h27186;
         mem[625] =  20'h3410a;
         mem[626] =  20'h1ac90;
         mem[627] =  20'h34124;
         mem[628] =  20'h0ddc9;
         mem[629] =  20'h64e68;
         mem[630] =  20'h00148;
         mem[631] =  20'h0de12;
         mem[632] =  20'h44f0b;
         mem[633] =  20'h13a45;
         mem[634] =  20'h64643;
         mem[635] =  20'h6ba43;
         mem[636] =  20'h51926;
         mem[637] =  20'h38aea;
         mem[638] =  20'h2ca43;
         mem[639] =  20'h33983;
         mem[640] =  20'h0e076;
         mem[641] =  20'h6dd46;
         mem[642] =  20'h70d46;
         mem[643] =  20'h158cc;
         mem[644] =  20'h28089;
         mem[645] =  20'h02cc9;
         mem[646] =  20'h01cc9;
         mem[647] =  20'h41926;
         mem[648] =  20'h454c9;
         mem[649] =  20'h22c73;
         mem[650] =  20'h27126;
         mem[651] =  20'h22c73;
         mem[652] =  20'h12cc9;
         mem[653] =  20'h84a43;
         mem[654] =  20'h3ee44;
         mem[655] =  20'h1c50a;
         mem[656] =  20'h33d26;
         mem[657] =  20'h3b528;
         mem[658] =  20'h258ac;
         mem[659] =  20'h275c6;
         mem[660] =  20'h21073;
         mem[661] =  20'h1b1f4;
         mem[662] =  20'h195f4;
         mem[663] =  20'h41cc6;
         mem[664] =  20'h3fcc6;
         mem[665] =  20'h100ce;
         mem[666] =  20'h0d8ce;
         mem[667] =  20'h1c0c7;
         mem[668] =  20'h1b4c9;
         mem[669] =  20'h1bd0a;
         mem[670] =  20'h1a50a;
         mem[671] =  20'h72946;
         mem[672] =  20'h70ea6;
         mem[673] =  20'h0ed86;
         mem[674] =  20'h0d586;
         mem[675] =  20'h22586;
         mem[676] =  20'h340c9;
         mem[677] =  20'h2c686;
         mem[678] =  20'h1f586;
         mem[679] =  20'h5b10a;
         mem[680] =  20'h5810a;
         mem[681] =  20'h4568d;
         mem[682] =  20'h39d85;
         mem[683] =  20'h26e06;
         mem[684] =  20'h77124;
         mem[685] =  20'h21185;
         mem[686] =  20'h201cc;
         mem[687] =  20'h1b526;
         mem[688] =  20'h26263;
         mem[689] =  20'h430c9;
         mem[690] =  20'h2ca42;
         mem[691] =  20'h11892;
         mem[692] =  20'h71283;
         mem[693] =  20'h38ac3;
         mem[694] =  20'h0c892;
         mem[695] =  20'h04c97;
         mem[696] =  20'h12cd3;
         mem[697] =  20'h110c9;
         mem[698] =  20'h1f546;
         mem[699] =  20'h01d8c;
         mem[700] =  20'h12f06;
         mem[701] =  20'h5a08a;
         mem[702] =  20'h3a48f;
         mem[703] =  20'h45e26;
         mem[704] =  20'h1fe48;
         mem[705] =  20'h275c6;
         mem[706] =  20'h265c6;
         mem[707] =  20'h23472;
         mem[708] =  20'h20872;
         mem[709] =  20'h411c4;
         mem[710] =  20'h3f924;
         mem[711] =  20'h00a49;
         mem[712] =  20'h14588;
         mem[713] =  20'h06905;
         mem[714] =  20'h2ece8;
         mem[715] =  20'h4b2c4;
         mem[716] =  20'h2948f;
         mem[717] =  20'h2d0e8;
         mem[718] =  20'h72924;
         mem[719] =  20'h0cec4;
         mem[720] =  20'h170d1;
         mem[721] =  20'h0e912;
         mem[722] =  20'h044cc;
         mem[723] =  20'h01cc9;
         mem[724] =  20'h2312c;
         mem[725] =  20'h8a242;
         mem[726] =  20'h41186;
         mem[727] =  20'h0648b;
         mem[728] =  20'h0508a;
         mem[729] =  20'h130d1;
         mem[730] =  20'h61926;
         mem[731] =  20'h51509;
         mem[732] =  20'h360cc;
         mem[733] =  20'h328cc;
         mem[734] =  20'h0f08f;
         mem[735] =  20'h1fa63;
         mem[736] =  20'h34d27;
         mem[737] =  20'h32d89;
         mem[738] =  20'h26643;
         mem[739] =  20'h0288c;
         mem[740] =  20'h3924e;
         mem[741] =  20'h00089;
         mem[742] =  20'h22492;
         mem[743] =  20'h21492;
         mem[744] =  20'h21cca;
         mem[745] =  20'h1b48b;
         mem[746] =  20'h65243;
         mem[747] =  20'h64283;
         mem[748] =  20'h3a8cc;
         mem[749] =  20'h53508;
         mem[750] =  20'h41c6c;
         mem[751] =  20'h399ce;
         mem[752] =  20'h0030a;
         mem[753] =  20'h45242;
         mem[754] =  20'h240ac;
         mem[755] =  20'h1f4ac;
         mem[756] =  20'h29912;
         mem[757] =  20'h25912;
         mem[758] =  20'h2258c;
         mem[759] =  20'h274c9;
         mem[760] =  20'h538cb;
         mem[761] =  20'h1f58c;
         mem[762] =  20'h0cee3;
         mem[763] =  20'h5e263;
         mem[764] =  20'h6d964;
         mem[765] =  20'h51505;
         mem[766] =  20'h41944;
         mem[767] =  20'h26929;
         mem[768] =  20'h5b526;
         mem[769] =  20'h4b526;
         mem[770] =  20'h3f688;
         mem[771] =  20'h00932;
         mem[772] =  20'h4812a;
         mem[773] =  20'h0cd05;
         mem[774] =  20'h19ea6;
         mem[775] =  20'h01d4e;
         mem[776] =  20'h6d584;
         mem[777] =  20'h25ae4;
         mem[778] =  20'h41d0a;
         mem[779] =  20'h64243;
         mem[780] =  20'h67d24;
         mem[781] =  20'h64124;
         mem[782] =  20'h480c6;
         mem[783] =  20'h460c6;
         mem[784] =  20'h12f06;
         mem[785] =  20'h19a43;
         mem[786] =  20'h00304;
         mem[787] =  20'h64643;
         mem[788] =  20'h61926;
         mem[789] =  20'h5dd26;
         mem[790] =  20'h6be43;
         mem[791] =  20'h340ca;
         mem[792] =  20'h280c9;
         mem[793] =  20'h340a8;
         mem[794] =  20'h350c8;
         mem[795] =  20'h20ccb;
         mem[796] =  20'h28d09;
         mem[797] =  20'h2c2a6;
         mem[798] =  20'h2306c;
         mem[799] =  20'h39d6c;
         mem[800] =  20'h35548;
         mem[801] =  20'h33583;
         mem[802] =  20'h46644;
         mem[803] =  20'h002d6;
         mem[804] =  20'h0f4c8;
         mem[805] =  20'h024c9;
         mem[806] =  20'h028c9;
         mem[807] =  20'h14cce;
         mem[808] =  20'h3f648;
         mem[809] =  20'h0286e;
         mem[810] =  20'h13e14;
         mem[811] =  20'h1b4ca;
         mem[812] =  20'h01604;
         mem[813] =  20'h1fe44;
         mem[814] =  20'h034c9;
         mem[815] =  20'h1b105;
         mem[816] =  20'h41944;
         mem[817] =  20'h3f144;
         mem[818] =  20'h46985;
         mem[819] =  20'h3f50a;
         mem[820] =  20'h4dd28;
         mem[821] =  20'h83703;
         mem[822] =  20'h7de44;
         mem[823] =  20'h5e126;
         mem[824] =  20'h6d144;
         mem[825] =  20'h4d48c;
         mem[826] =  20'h27d26;
         mem[827] =  20'h518c9;
         mem[828] =  20'h65984;
         mem[829] =  20'h1fa83;
         mem[830] =  20'h08529;
         mem[831] =  20'h77524;
         mem[832] =  20'h09092;
         mem[833] =  20'h0e50c;
         mem[834] =  20'h41528;
         mem[835] =  20'h46185;
         mem[836] =  20'h3b126;
         mem[837] =  20'h3fcc9;
         mem[838] =  20'h2ccac;
         mem[839] =  20'h00aa6;
         mem[840] =  20'h27546;
         mem[841] =  20'h024cf;
         mem[842] =  20'h0d242;
         mem[843] =  20'h6c506;
         mem[844] =  20'h00e42;
         mem[845] =  20'h02126;
         mem[846] =  20'h6a643;
         mem[847] =  20'h2d585;
         mem[848] =  20'h12cc9;
         mem[849] =  20'h11889;
         mem[850] =  20'h0c889;
         mem[851] =  20'h06704;
         mem[852] =  20'h64126;
         mem[853] =  20'h54d26;
         mem[854] =  20'h5de63;
         mem[855] =  20'h1facc;
         mem[856] =  20'h528c6;
         mem[857] =  20'h0da83;
         mem[858] =  20'h598ca;
         mem[859] =  20'h4ca06;
         mem[860] =  20'h51d09;
         mem[861] =  20'h34cce;
         mem[862] =  20'h4ba06;
         mem[863] =  20'h65608;
         mem[864] =  20'h0888c;
         mem[865] =  20'h0e90a;
         mem[866] =  20'h27186;
         mem[867] =  20'h2e4c9;
         mem[868] =  20'h0010c;
         mem[869] =  20'h368c9;
         mem[870] =  20'h4b8c6;
         mem[871] =  20'h842a3;
         mem[872] =  20'h00a06;
         mem[873] =  20'h28ce6;
         mem[874] =  20'h1a88e;
         mem[875] =  20'h2e0c9;
         mem[876] =  20'h33cce;
         mem[877] =  20'h36890;
         mem[878] =  20'h59cca;
         mem[879] =  20'h46585;
         mem[880] =  20'h4b2e3;
         mem[881] =  20'h034cc;
         mem[882] =  20'h3e985;
         mem[883] =  20'h0fd44;
         mem[884] =  20'h014cc;
         mem[885] =  20'h28526;
         mem[886] =  20'h26926;
         mem[887] =  20'h4664d;
         mem[888] =  20'h44e4d;
         mem[889] =  20'h67186;
         mem[890] =  20'h25aa3;
         mem[891] =  20'h67186;
         mem[892] =  20'h2d0ce;
         mem[893] =  20'h3fe62;
         mem[894] =  20'h1a5c4;
         mem[895] =  20'h71644;
         mem[896] =  20'h01c89;
         mem[897] =  20'h16164;
         mem[898] =  20'h00926;
         mem[899] =  20'h0b097;
         mem[900] =  20'h06897;
         mem[901] =  20'h65643;
         mem[902] =  20'h12d64;
         mem[903] =  20'h64a83;
         mem[904] =  20'h141a4;
         mem[905] =  20'h38acf;
         mem[906] =  20'h19dc3;
         mem[907] =  20'h2dd44;
         mem[908] =  20'h2d544;
         mem[909] =  20'h1b8c9;
         mem[910] =  20'h4b526;
         mem[911] =  20'h14d0a;
         mem[912] =  20'h26606;
         mem[913] =  20'h26dc6;
         mem[914] =  20'h13d26;
         mem[915] =  20'h14642;
         mem[916] =  20'h27526;
         mem[917] =  20'h06703;
         mem[918] =  20'h6a546;
         mem[919] =  20'h71643;
         mem[920] =  20'h1fcd0;
         mem[921] =  20'h27566;
         mem[922] =  20'h0dd96;
         mem[923] =  20'h2e48a;
         mem[924] =  20'h02492;
         mem[925] =  20'h368c9;
         mem[926] =  20'h2cdea;
         mem[927] =  20'h21cc9;
         mem[928] =  20'h3a8ca;
         mem[929] =  20'h5a4ca;
         mem[930] =  20'h594ca;
         mem[931] =  20'h33209;
         mem[932] =  20'h45683;
         mem[933] =  20'h0348d;
         mem[934] =  20'h01c8d;
         mem[935] =  20'h07247;
         mem[936] =  20'h450c9;
         mem[937] =  20'h72926;
         mem[938] =  20'h391e6;
         mem[939] =  20'h3fe62;
         mem[940] =  20'h278f0;
         mem[941] =  20'h59d26;
         mem[942] =  20'h2bd0c;
         mem[943] =  20'h1aa43;
         mem[944] =  20'h64186;
         mem[945] =  20'h54924;
         mem[946] =  20'h335ce;
         mem[947] =  20'h646c6;
         mem[948] =  20'h024c9;
         mem[949] =  20'h2194a;
         mem[950] =  20'h2094a;
         mem[951] =  20'h26a06;
         mem[952] =  20'h2bcc9;
         mem[953] =  20'h4290e;
         mem[954] =  20'h4d4cc;
         mem[955] =  20'h4090c;
         mem[956] =  20'h02089;
         mem[957] =  20'h1b910;
         mem[958] =  20'h40546;
         mem[959] =  20'h26dce;
         mem[960] =  20'h45682;
         mem[961] =  20'h36890;
         mem[962] =  20'h4518a;
         mem[963] =  20'h39d84;
         mem[964] =  20'h4d4c7;
         mem[965] =  20'h1b910;
         mem[966] =  20'h1a910;
         mem[967] =  20'h3a526;
         mem[968] =  20'h1fa0c;
         mem[969] =  20'h3a8c8;
         mem[970] =  20'h01872;
         mem[971] =  20'h3c8ae;
         mem[972] =  20'h38cae;
         mem[973] =  20'h1ad46;
         mem[974] =  20'h132f2;
         mem[975] =  20'h06aa3;
         mem[976] =  20'h27cc9;
         mem[977] =  20'h71586;
         mem[978] =  20'h36110;
         mem[979] =  20'h76f04;
         mem[980] =  20'h36110;
         mem[981] =  20'h32110;
         mem[982] =  20'h4d10a;
         mem[983] =  20'h2d0a8;
         mem[984] =  20'h07662;
         mem[985] =  20'h4b309;
         mem[986] =  20'h019a8;
         mem[987] =  20'h00303;
         mem[988] =  20'h17c8b;
         mem[989] =  20'h278c9;
         mem[990] =  20'h46588;
         mem[991] =  20'h32186;
         mem[992] =  20'h6be43;
         mem[993] =  20'h57926;
         mem[994] =  20'h17c89;
         mem[995] =  20'h12c89;
         mem[996] =  20'h03d33;
         mem[997] =  20'h00133;
         mem[998] =  20'h480c8;
         mem[999] =  20'h460c8;
         mem[1000] =  20'h46263;
         mem[1001] =  20'h7de44;
         mem[1002] =  20'h27206;
         mem[1003] =  20'h01926;
         mem[1004] =  20'h1548e;
         mem[1005] =  20'h1f9ec;
         mem[1006] =  20'h4dd05;
         mem[1007] =  20'h014c9;
         mem[1008] =  20'h030c9;
         mem[1009] =  20'h20988;
         mem[1010] =  20'h4e566;
         mem[1011] =  20'h516a3;
         mem[1012] =  20'h0850c;
         mem[1013] =  20'h004cc;
         mem[1014] =  20'h0d2a2;
         mem[1015] =  20'h0d263;
         mem[1016] =  20'h42cce;
         mem[1017] =  20'h3ecce;
         mem[1018] =  20'h275ce;
         mem[1019] =  20'h4b126;
         mem[1020] =  20'h5b509;
         mem[1021] =  20'h06ac4;
         mem[1022] =  20'h47126;
         mem[1023] =  20'h5de43;
         mem[1024] =  20'h5b8e9;
         mem[1025] =  20'h13e04;
         mem[1026] =  20'h27585;
         mem[1027] =  20'h27c89;
         mem[1028] =  20'h0948a;
         mem[1029] =  20'h0848a;
         mem[1030] =  20'h618c9;
         mem[1031] =  20'h5e8c9;
         mem[1032] =  20'h0a073;
         mem[1033] =  20'h130c9;
         mem[1034] =  20'h03c73;
         mem[1035] =  20'h14584;
         mem[1036] =  20'h21c89;
         mem[1037] =  20'h01873;
         mem[1038] =  20'h0906c;
         mem[1039] =  20'h2d545;
         mem[1040] =  20'h15872;
         mem[1041] =  20'h150cc;
         mem[1042] =  20'h2ca63;
         mem[1043] =  20'h2c643;
         mem[1044] =  20'h52244;
         mem[1045] =  20'h200c9;
         mem[1046] =  20'h07684;
         mem[1047] =  20'h06684;
         mem[1048] =  20'h604c6;
         mem[1049] =  20'h0cb08;
         mem[1050] =  20'h20a43;
         mem[1051] =  20'h5fcc6;
         mem[1052] =  20'h4dd05;
         mem[1053] =  20'h4c505;
         mem[1054] =  20'h015c6;
         mem[1055] =  20'h0f08f;
         mem[1056] =  20'h2e4ac;
         mem[1057] =  20'h3a10e;
         mem[1058] =  20'h1fac6;
         mem[1059] =  20'h1f4c6;
         mem[1060] =  20'h6d524;
         mem[1061] =  20'h71263;
         mem[1062] =  20'h6d524;
         mem[1063] =  20'h6aa43;
         mem[1064] =  20'h6d524;
         mem[1065] =  20'h00303;
         mem[1066] =  20'h015c4;
         mem[1067] =  20'h59126;
         mem[1068] =  20'h54cc9;
         mem[1069] =  20'h7e5a4;
         mem[1070] =  20'h3a8cc;
         mem[1071] =  20'h3eea3;
         mem[1072] =  20'h34126;
         mem[1073] =  20'h3f527;
         mem[1074] =  20'h41948;
         mem[1075] =  20'h5df03;
         mem[1076] =  20'h21526;
         mem[1077] =  20'h524c9;
         mem[1078] =  20'h6d524;
         mem[1079] =  20'h4d4c6;
         mem[1080] =  20'h3a9ca;
         mem[1081] =  20'h389ca;
         mem[1082] =  20'h2dd31;
         mem[1083] =  20'h19cd4;
         mem[1084] =  20'h33d44;
         mem[1085] =  20'h2e489;
         mem[1086] =  20'h604c9;
         mem[1087] =  20'h32cd0;
         mem[1088] =  20'h6d524;
         mem[1089] =  20'h6b124;
         mem[1090] =  20'h08d26;
         mem[1091] =  20'h2d08a;
         mem[1092] =  20'h21186;
         mem[1093] =  20'h1a928;
         mem[1094] =  20'h67148;
         mem[1095] =  20'h64948;
         mem[1096] =  20'h00304;
         mem[1097] =  20'h25926;
         mem[1098] =  20'h19306;
         mem[1099] =  20'h01564;
         mem[1100] =  20'h06ac4;
         mem[1101] =  20'h27cd2;
         mem[1102] =  20'h38e84;
         mem[1103] =  20'h0ddce;
         mem[1104] =  20'h0da06;
         mem[1105] =  20'h13663;
         mem[1106] =  20'h08144;
         mem[1107] =  20'h3848f;
         mem[1108] =  20'h3f2a3;
         mem[1109] =  20'h00cc6;
         mem[1110] =  20'h1a9c9;
         mem[1111] =  20'h088c9;
         mem[1112] =  20'h35d29;
         mem[1113] =  20'h02095;
         mem[1114] =  20'h8a662;
         mem[1115] =  20'h5e683;
         mem[1116] =  20'h04c8d;
         mem[1117] =  20'h2c108;
         mem[1118] =  20'h5b0c9;
         mem[1119] =  20'h588c9;
         mem[1120] =  20'h22c8a;
         mem[1121] =  20'h20c8a;
         mem[1122] =  20'h22cc6;
         mem[1123] =  20'h204c6;
         mem[1124] =  20'h0cb15;
         mem[1125] =  20'h0cccd;
         mem[1126] =  20'h05095;
         mem[1127] =  20'h19094;
         mem[1128] =  20'h66126;
         mem[1129] =  20'h01cc9;
         mem[1130] =  20'h4f0e9;
         mem[1131] =  20'h849c3;
         mem[1132] =  20'h220c9;
         mem[1133] =  20'h21c8a;
         mem[1134] =  20'h280c9;
         mem[1135] =  20'h210c9;
         mem[1136] =  20'h5b144;
         mem[1137] =  20'h209ce;
         mem[1138] =  20'h35186;
         mem[1139] =  20'h2718c;
         mem[1140] =  20'h540ca;
         mem[1141] =  20'h3ee88;
         mem[1142] =  20'h55126;
         mem[1143] =  20'h024c9;
         mem[1144] =  20'h08cae;
         mem[1145] =  20'h19e06;
         mem[1146] =  20'h16d09;
         mem[1147] =  20'h530ca;
         mem[1148] =  20'h55126;
         mem[1149] =  20'h51526;
         mem[1150] =  20'h67526;
         mem[1151] =  20'h64926;
         mem[1152] =  20'h65643;
         mem[1153] =  20'h64643;
         mem[1154] =  20'h01643;
         mem[1155] =  20'h06a62;
         mem[1156] =  20'h100cb;
         mem[1157] =  20'h5ede6;
         mem[1158] =  20'h100cb;
         mem[1159] =  20'h0d8cb;
         mem[1160] =  20'h110c9;
         mem[1161] =  20'h0cec4;
         mem[1162] =  20'h00aac;
         mem[1163] =  20'h4b243;
         mem[1164] =  20'h0f8c9;
         mem[1165] =  20'h3f643;
         mem[1166] =  20'h16d09;
         mem[1167] =  20'h2ca43;
         mem[1168] =  20'h470c9;
         mem[1169] =  20'h344c9;
         mem[1170] =  20'h03c52;
         mem[1171] =  20'h01c52;
         mem[1172] =  20'h170e9;
         mem[1173] =  20'h71526;
         mem[1174] =  20'h716a3;
         mem[1175] =  20'h12ce9;
         mem[1176] =  20'h2c6c3;
         mem[1177] =  20'h12f10;
         mem[1178] =  20'h6d924;
         mem[1179] =  20'h20988;
         mem[1180] =  20'h26dc6;
         mem[1181] =  20'h655c6;
         mem[1182] =  20'h110c9;
         mem[1183] =  20'h0c8c9;
         mem[1184] =  20'h19e8a;
         mem[1185] =  20'h51d28;
         mem[1186] =  20'h06eaf;
         mem[1187] =  20'h4c5c8;
         mem[1188] =  20'h2d584;
         mem[1189] =  20'h20d26;
         mem[1190] =  20'h480c6;
         mem[1191] =  20'h460c6;
         mem[1192] =  20'h1aa42;
         mem[1193] =  20'h0c8cb;
         mem[1194] =  20'h048cf;
         mem[1195] =  20'h000cd;
         mem[1196] =  20'h030c9;
         mem[1197] =  20'h018c9;
         mem[1198] =  20'h0cb04;
         mem[1199] =  20'h52244;
         mem[1200] =  20'h2e144;
         mem[1201] =  20'h33583;
         mem[1202] =  20'h58a63;
         mem[1203] =  20'h02894;
         mem[1204] =  20'h5fd26;
         mem[1205] =  20'h38de4;
         mem[1206] =  20'h1b187;
         mem[1207] =  20'h3e8c9;
         mem[1208] =  20'h23cc9;
         mem[1209] =  20'h70a06;
         mem[1210] =  20'h72dc6;
         mem[1211] =  20'h7d684;
         mem[1212] =  20'h32a86;
         mem[1213] =  20'h33cc9;
         mem[1214] =  20'h21588;
         mem[1215] =  20'h20588;
         mem[1216] =  20'h280c9;
         mem[1217] =  20'h008d0;
         mem[1218] =  20'h1cccc;
         mem[1219] =  20'h19ccc;
         mem[1220] =  20'h4ed26;
         mem[1221] =  20'h011f6;
         mem[1222] =  20'h4ed26;
         mem[1223] =  20'h4b126;
         mem[1224] =  20'h61926;
         mem[1225] =  20'h5dd26;
         mem[1226] =  20'h0290a;
         mem[1227] =  20'h00490;
         mem[1228] =  20'h27546;
         mem[1229] =  20'h4d88a;
         mem[1230] =  20'h1b146;
         mem[1231] =  20'h8a642;
         mem[1232] =  20'h2d966;
         mem[1233] =  20'h0018a;
         mem[1234] =  20'h08d86;
         mem[1235] =  20'h65d24;
         mem[1236] =  20'h2d1f0;
         mem[1237] =  20'h3fd8d;
         mem[1238] =  20'h0e186;
         mem[1239] =  20'h39189;
         mem[1240] =  20'h10906;
         mem[1241] =  20'h0c906;
         mem[1242] =  20'h12f0b;
         mem[1243] =  20'h5150a;
         mem[1244] =  20'h5a08a;
         mem[1245] =  20'h0f095;
         mem[1246] =  20'h1a1e9;
         mem[1247] =  20'h06706;
         mem[1248] =  20'h27cb0;
         mem[1249] =  20'h84243;
         mem[1250] =  20'h20c6c;
         mem[1251] =  20'h28489;
         mem[1252] =  20'h26d28;
         mem[1253] =  20'h13e82;
         mem[1254] =  20'h3f243;
         mem[1255] =  20'h5f946;
         mem[1256] =  20'h19492;
         mem[1257] =  20'h034c9;
         mem[1258] =  20'h014c9;
         mem[1259] =  20'h02cc9;
         mem[1260] =  20'h2d526;
         mem[1261] =  20'h00e42;
         mem[1262] =  20'h3ea84;
         mem[1263] =  20'h0f08c;
         mem[1264] =  20'h20ccc;
         mem[1265] =  20'h01a56;
         mem[1266] =  20'h00256;
         mem[1267] =  20'h110cb;
         mem[1268] =  20'h0c8cb;
         mem[1269] =  20'h02cc9;
         mem[1270] =  20'h00283;
         mem[1271] =  20'h0d282;
         mem[1272] =  20'h3ee42;
         mem[1273] =  20'h304c9;
         mem[1274] =  20'h002c9;
         mem[1275] =  20'h170c9;
         mem[1276] =  20'h2bcc9;
         mem[1277] =  20'h25b06;
         mem[1278] =  20'h0c8ca;
         mem[1279] =  20'h280c9;
         mem[1280] =  20'h01cc9;
         mem[1281] =  20'h03cc9;
         mem[1282] =  20'h00cc9;
         mem[1283] =  20'h6e126;
         mem[1284] =  20'h6a643;
         mem[1285] =  20'h5b526;
         mem[1286] =  20'h5dee6;
         mem[1287] =  20'h5f243;
         mem[1288] =  20'h57926;
         mem[1289] =  20'h3450a;
         mem[1290] =  20'h2c9e6;
         mem[1291] =  20'h3450a;
         mem[1292] =  20'h014cc;
         mem[1293] =  20'h3450a;
         mem[1294] =  20'h214c9;
         mem[1295] =  20'h28092;
         mem[1296] =  20'h2d184;
         mem[1297] =  20'h3450a;
         mem[1298] =  20'h33d0a;
         mem[1299] =  20'h414ce;
         mem[1300] =  20'h218d3;
         mem[1301] =  20'h4c986;
         mem[1302] =  20'h38a46;
         mem[1303] =  20'h5b90a;
         mem[1304] =  20'h386c8;
         mem[1305] =  20'h72986;
         mem[1306] =  20'h25a92;
         mem[1307] =  20'h2668c;
         mem[1308] =  20'h64148;
         mem[1309] =  20'h65a43;
         mem[1310] =  20'h44e63;
         mem[1311] =  20'h290c9;
         mem[1312] =  20'h2c2c4;
         mem[1313] =  20'h28cec;
         mem[1314] =  20'h2cd69;
         mem[1315] =  20'h41948;
         mem[1316] =  20'h4b927;
         mem[1317] =  20'h5b8c9;
         mem[1318] =  20'h4bccc;
         mem[1319] =  20'h54cc6;
         mem[1320] =  20'h020c9;
         mem[1321] =  20'h088d7;
         mem[1322] =  20'h64126;
         mem[1323] =  20'h6b643;
         mem[1324] =  20'h0ddae;
         mem[1325] =  20'h03d0c;
         mem[1326] =  20'h0010c;
         mem[1327] =  20'h0e907;
         mem[1328] =  20'h068c9;
         mem[1329] =  20'h358cc;
         mem[1330] =  20'h330cc;
         mem[1331] =  20'h234af;
         mem[1332] =  20'h200af;
         mem[1333] =  20'h1d8c9;
         mem[1334] =  20'h2c0cf;
         mem[1335] =  20'h60988;
         mem[1336] =  20'h0cb04;
         mem[1337] =  20'h0a053;
         mem[1338] =  20'h08053;
         mem[1339] =  20'h0bc54;
         mem[1340] =  20'h06454;
         mem[1341] =  20'h494cc;
         mem[1342] =  20'h44ccc;
         mem[1343] =  20'h2664e;
         mem[1344] =  20'h400e8;
         mem[1345] =  20'h3a18c;
         mem[1346] =  20'h71245;
         mem[1347] =  20'h84683;
         mem[1348] =  20'h4d4cc;
         mem[1349] =  20'h26a43;
         mem[1350] =  20'h26643;
         mem[1351] =  20'h1d8c9;
         mem[1352] =  20'h4b926;
         mem[1353] =  20'h58a44;
         mem[1354] =  20'h2d8ce;
         mem[1355] =  20'h53186;
         mem[1356] =  20'h2d589;
         mem[1357] =  20'h4e0c6;
         mem[1358] =  20'h0c88a;
         mem[1359] =  20'h02126;
         mem[1360] =  20'h38d86;
         mem[1361] =  20'h41cc9;
         mem[1362] =  20'h3fcc9;
         mem[1363] =  20'h60126;
         mem[1364] =  20'h65586;
         mem[1365] =  20'h0d683;
         mem[1366] =  20'h1fd86;
         mem[1367] =  20'h02c78;
         mem[1368] =  20'h64de4;
         mem[1369] =  20'h4d4cc;
         mem[1370] =  20'h5e188;
         mem[1371] =  20'h4250e;
         mem[1372] =  20'h3890e;
         mem[1373] =  20'h4712a;
         mem[1374] =  20'h2d586;
         mem[1375] =  20'h604c9;
         mem[1376] =  20'h33d27;
         mem[1377] =  20'h1b90a;
         mem[1378] =  20'h268c9;
         mem[1379] =  20'h25b0c;
         mem[1380] =  20'h2c8ce;
         mem[1381] =  20'h36ca8;
         mem[1382] =  20'h320a8;
         mem[1383] =  20'h170c6;
         mem[1384] =  20'h130c6;
         mem[1385] =  20'h110c9;
         mem[1386] =  20'h0c8c9;
         mem[1387] =  20'h13a46;
         mem[1388] =  20'h13526;
         mem[1389] =  20'h15148;
         mem[1390] =  20'h14148;
         mem[1391] =  20'h474cc;
         mem[1392] =  20'h46ccb;
         mem[1393] =  20'h33d44;
         mem[1394] =  20'h27cc7;
         mem[1395] =  20'h71e43;
         mem[1396] =  20'h1b0c9;
         mem[1397] =  20'h08527;
         mem[1398] =  20'h464c6;
         mem[1399] =  20'h4e88b;
         mem[1400] =  20'h4c88b;
         mem[1401] =  20'h02192;
         mem[1402] =  20'h4b945;
         mem[1403] =  20'h7dac3;
         mem[1404] =  20'h19054;
         mem[1405] =  20'h0cb04;
         mem[1406] =  20'h33d44;
         mem[1407] =  20'h2d50a;
         mem[1408] =  20'h038ce;
         mem[1409] =  20'h45ca8;
         mem[1410] =  20'h00a89;
         mem[1411] =  20'h2d588;
         mem[1412] =  20'h6c8c6;
         mem[1413] =  20'h40544;
         mem[1414] =  20'h20d89;
         mem[1415] =  20'h460c8;
         mem[1416] =  20'h1d891;
         mem[1417] =  20'h000c6;
         mem[1418] =  20'h1d891;
         mem[1419] =  20'h19891;
         mem[1420] =  20'h71e63;
         mem[1421] =  20'h02c52;
         mem[1422] =  20'h1cc52;
         mem[1423] =  20'h1ac52;
         mem[1424] =  20'h46948;
         mem[1425] =  20'h28089;
         mem[1426] =  20'h028c9;
         mem[1427] =  20'h38e08;
         mem[1428] =  20'h614c9;
         mem[1429] =  20'h2dcc9;
         mem[1430] =  20'h614c9;
         mem[1431] =  20'h4bd86;
         mem[1432] =  20'h4e926;
         mem[1433] =  20'h4b526;
         mem[1434] =  20'h2ca43;
         mem[1435] =  20'h2c2c6;
         mem[1436] =  20'h1d8c6;
         mem[1437] =  20'h190c6;
         mem[1438] =  20'h46206;
         mem[1439] =  20'h65924;
         mem[1440] =  20'h614c9;
         mem[1441] =  20'h5ecc9;
         mem[1442] =  20'h0a0d7;
         mem[1443] =  20'h83703;
         mem[1444] =  20'h7d304;
         mem[1445] =  20'h070d7;
         mem[1446] =  20'h6b243;
         mem[1447] =  20'h64243;
         mem[1448] =  20'h646c4;
         mem[1449] =  20'h64126;
         mem[1450] =  20'h3f2a3;
         mem[1451] =  20'h71186;
         mem[1452] =  20'h1f704;
         mem[1453] =  20'h0f08f;
         mem[1454] =  20'h2e4cc;
         mem[1455] =  20'h270c9;
         mem[1456] =  20'h02cc9;
         mem[1457] =  20'h2e0c9;
         mem[1458] =  20'h06e83;
         mem[1459] =  20'h70d86;
         mem[1460] =  20'h0fc8d;
         mem[1461] =  20'h2d584;
         mem[1462] =  20'h08c8d;
         mem[1463] =  20'h01872;
         mem[1464] =  20'h16545;
         mem[1465] =  20'h5f588;
         mem[1466] =  20'h40cc9;
         mem[1467] =  20'h14c89;
         mem[1468] =  20'h044ce;
         mem[1469] =  20'h004ce;
         mem[1470] =  20'h038d0;
         mem[1471] =  20'h1ac8a;
         mem[1472] =  20'h6b246;
         mem[1473] =  20'h7d6c4;
         mem[1474] =  20'h16545;
         mem[1475] =  20'h12d45;
         mem[1476] =  20'h28990;
         mem[1477] =  20'h25990;
         mem[1478] =  20'h3acaf;
         mem[1479] =  20'h70ea2;
         mem[1480] =  20'h03d26;
         mem[1481] =  20'h07d84;
         mem[1482] =  20'h0198c;
         mem[1483] =  20'h4090c;
         mem[1484] =  20'h67948;
         mem[1485] =  20'h64148;
         mem[1486] =  20'h4d985;
         mem[1487] =  20'h65948;
         mem[1488] =  20'h27586;
         mem[1489] =  20'h27c92;
         mem[1490] =  20'h3acce;
         mem[1491] =  20'h3a4ce;
         mem[1492] =  20'h1ad6c;
         mem[1493] =  20'h330d0;
         mem[1494] =  20'h17095;
         mem[1495] =  20'h13895;
         mem[1496] =  20'h08d12;
         mem[1497] =  20'h1fe08;
         mem[1498] =  20'h2664c;
         mem[1499] =  20'h3fa0c;
         mem[1500] =  20'h1cd14;
         mem[1501] =  20'h0e526;
         mem[1502] =  20'h1cd14;
         mem[1503] =  20'h19514;
         mem[1504] =  20'h34d0e;
         mem[1505] =  20'h3350e;
         mem[1506] =  20'h53ca8;
         mem[1507] =  20'h524e9;
         mem[1508] =  20'h5170a;
         mem[1509] =  20'h0d90b;
         mem[1510] =  20'h0f110;
         mem[1511] =  20'h0cb06;
         mem[1512] =  20'h01989;
         mem[1513] =  20'h0cd8c;
         mem[1514] =  20'h23cc9;
         mem[1515] =  20'h13d0a;
         mem[1516] =  20'h84e43;
         mem[1517] =  20'h3ee42;
         mem[1518] =  20'h3eec3;
         mem[1519] =  20'h32989;
         mem[1520] =  20'h35186;
         mem[1521] =  20'h32186;
         mem[1522] =  20'h604c9;
         mem[1523] =  20'h53126;
         mem[1524] =  20'h344ec;
         mem[1525] =  20'h52526;
         mem[1526] =  20'h5f644;
         mem[1527] =  20'h1a490;
         mem[1528] =  20'h604c9;
         mem[1529] =  20'h5fcc9;
         mem[1530] =  20'h4718a;
         mem[1531] =  20'h265c6;
         mem[1532] =  20'h0da28;
         mem[1533] =  20'h0e195;
         mem[1534] =  20'h08529;
         mem[1535] =  20'h2bf03;
         mem[1536] =  20'h2852a;
         mem[1537] =  20'h45643;
         mem[1538] =  20'h66124;
         mem[1539] =  20'h00126;
         mem[1540] =  20'h44f06;
         mem[1541] =  20'h38e86;
         mem[1542] =  20'h2060c;
         mem[1543] =  20'h0f08f;
         mem[1544] =  20'h14944;
         mem[1545] =  20'h600c8;
         mem[1546] =  20'h044ea;
         mem[1547] =  20'h000ea;
         mem[1548] =  20'h0a4cc;
         mem[1549] =  20'h00668;
         mem[1550] =  20'h0f924;
         mem[1551] =  20'h0d524;
         mem[1552] =  20'h0f946;
         mem[1553] =  20'h19e42;
         mem[1554] =  20'h09489;
         mem[1555] =  20'h08489;
         mem[1556] =  20'h21d0a;
         mem[1557] =  20'h1a98d;
         mem[1558] =  20'h228c6;
         mem[1559] =  20'h1f983;
         mem[1560] =  20'h21146;
         mem[1561] =  20'h00aa5;
         mem[1562] =  20'h32129;
         mem[1563] =  20'h27cc9;
         mem[1564] =  20'h12cc7;
         mem[1565] =  20'h72d86;
         mem[1566] =  20'h32a86;
         mem[1567] =  20'h0fd44;
         mem[1568] =  20'h204b2;
         mem[1569] =  20'h1e089;
         mem[1570] =  20'h2790e;
         mem[1571] =  20'h06706;
         mem[1572] =  20'h19089;
         mem[1573] =  20'h26643;
         mem[1574] =  20'h6b206;
         mem[1575] =  20'h28cc9;
         mem[1576] =  20'h26dc6;
         mem[1577] =  20'h2290a;
         mem[1578] =  20'h0d283;
         mem[1579] =  20'h0ed26;
         mem[1580] =  20'h278c9;
         mem[1581] =  20'h15c8b;
         mem[1582] =  20'h14c8b;
         mem[1583] =  20'h14d0a;
         mem[1584] =  20'h09052;
         mem[1585] =  20'h0ed26;
         mem[1586] =  20'h0ca63;
         mem[1587] =  20'h59d26;
         mem[1588] =  20'h32645;
         mem[1589] =  20'h030c9;
         mem[1590] =  20'h018c9;
         mem[1591] =  20'h28c8f;
         mem[1592] =  20'h1fa43;
         mem[1593] =  20'h2e1c6;
         mem[1594] =  20'h64a43;
         mem[1595] =  20'h6e126;
         mem[1596] =  20'h32186;
         mem[1597] =  20'h538e8;
         mem[1598] =  20'h6ae83;
         mem[1599] =  20'h6e126;
         mem[1600] =  20'h011e4;
         mem[1601] =  20'h10cc6;
         mem[1602] =  20'h12cc9;
         mem[1603] =  20'h6e126;
         mem[1604] =  20'h6a526;
         mem[1605] =  20'h72d86;
         mem[1606] =  20'h5e8c9;
         mem[1607] =  20'h5550a;
         mem[1608] =  20'h57b04;
         mem[1609] =  20'h73cc6;
         mem[1610] =  20'h5150a;
         mem[1611] =  20'h57b06;
         mem[1612] =  20'h0dd88;
         mem[1613] =  20'h3a526;
         mem[1614] =  20'h13e04;
         mem[1615] =  20'h0f08a;
         mem[1616] =  20'h1b0a8;
         mem[1617] =  20'h2212c;
         mem[1618] =  20'h2052c;
         mem[1619] =  20'h290c9;
         mem[1620] =  20'h19a8c;
         mem[1621] =  20'h1a230;
         mem[1622] =  20'h2dce6;
         mem[1623] =  20'h38ae2;
         mem[1624] =  20'h01cc9;
         mem[1625] =  20'h16089;
         mem[1626] =  20'h084cd;
         mem[1627] =  20'h8aa42;
         mem[1628] =  20'h3f526;
         mem[1629] =  20'h03858;
         mem[1630] =  20'h02058;
         mem[1631] =  20'h0d64a;
         mem[1632] =  20'h525e6;
         mem[1633] =  20'h84243;
         mem[1634] =  20'h0888b;
         mem[1635] =  20'h2e144;
         mem[1636] =  20'h01d52;
         mem[1637] =  20'h094d0;
         mem[1638] =  20'h07cd0;
         mem[1639] =  20'h110c6;
         mem[1640] =  20'h20242;
         mem[1641] =  20'h110c6;
         mem[1642] =  20'h0c8c6;
         mem[1643] =  20'h48166;
         mem[1644] =  20'h2d144;
         mem[1645] =  20'h3b147;
         mem[1646] =  20'h39147;
         mem[1647] =  20'h1d0c6;
         mem[1648] =  20'h26d48;
         mem[1649] =  20'h85203;
         mem[1650] =  20'h83a03;
         mem[1651] =  20'h1fece;
         mem[1652] =  20'h3f50a;
         mem[1653] =  20'h044cc;
         mem[1654] =  20'h0dcd2;
         mem[1655] =  20'h034c9;
         mem[1656] =  20'h4b0e9;
         mem[1657] =  20'h5510a;
         mem[1658] =  20'h004cc;
         mem[1659] =  20'h0946c;
         mem[1660] =  20'h5190a;
         mem[1661] =  20'h84262;
         mem[1662] =  20'h1448d;
         mem[1663] =  20'h3fe43;
         mem[1664] =  20'h150ac;
         mem[1665] =  20'h0f48f;
         mem[1666] =  20'h07604;
         mem[1667] =  20'h01a43;
         mem[1668] =  20'h07948;
         mem[1669] =  20'h73586;
         mem[1670] =  20'h5f183;
         mem[1671] =  20'h3eec4;
         mem[1672] =  20'h3a126;
         mem[1673] =  20'h46585;
         mem[1674] =  20'h2d547;
         mem[1675] =  20'h0f50a;
         mem[1676] =  20'h0dd0a;
         mem[1677] =  20'h1aa46;
         mem[1678] =  20'h1f549;
         mem[1679] =  20'h2c6a6;
         mem[1680] =  20'h192d0;
         mem[1681] =  20'h024d6;
         mem[1682] =  20'h0886c;
         mem[1683] =  20'h03192;
         mem[1684] =  20'h00192;
         mem[1685] =  20'h06ac4;
         mem[1686] =  20'h00e44;
         mem[1687] =  20'h1fec6;
         mem[1688] =  20'h014c9;
         mem[1689] =  20'h5a0c9;
         mem[1690] =  20'h598c9;
         mem[1691] =  20'h71e43;
         mem[1692] =  20'h018cd;
         mem[1693] =  20'h1ad84;
         mem[1694] =  20'h0dd86;
         mem[1695] =  20'h07643;
         mem[1696] =  20'h320cc;
         mem[1697] =  20'h600c9;
         mem[1698] =  20'h40ccd;
         mem[1699] =  20'h6be42;
         mem[1700] =  20'h1b4c9;
         mem[1701] =  20'h028c9;
         mem[1702] =  20'h26d48;
         mem[1703] =  20'h3bca8;
         mem[1704] =  20'h398a8;
         mem[1705] =  20'h48526;
         mem[1706] =  20'h0caef;
         mem[1707] =  20'h0410c;
         mem[1708] =  20'h5ecc9;
         mem[1709] =  20'h72924;
         mem[1710] =  20'h6a643;
         mem[1711] =  20'h48166;
         mem[1712] =  20'h44d66;
         mem[1713] =  20'h38706;
         mem[1714] =  20'h65908;
         mem[1715] =  20'h669c6;
         mem[1716] =  20'h06aa3;
         mem[1717] =  20'h0cb03;
         mem[1718] =  20'h5e505;
         mem[1719] =  20'h456a3;
         mem[1720] =  20'h70d86;
         mem[1721] =  20'h5a08a;
         mem[1722] =  20'h2d88a;
         mem[1723] =  20'h344cc;
         mem[1724] =  20'h08126;
         mem[1725] =  20'h58662;
         mem[1726] =  20'h2d94a;
         mem[1727] =  20'h4be4c;
         mem[1728] =  20'h020cc;
         mem[1729] =  20'h00e29;
         mem[1730] =  20'h0198b;
         mem[1731] =  20'h004cd;
         mem[1732] =  20'h33606;
         mem[1733] =  20'h340ac;
         mem[1734] =  20'h84243;
         mem[1735] =  20'h000c6;
         mem[1736] =  20'h00a83;
         mem[1737] =  20'h269ea;
         mem[1738] =  20'h27cc9;
         mem[1739] =  20'h024c9;
         mem[1740] =  20'h038c9;
         mem[1741] =  20'h65d26;
         mem[1742] =  20'h038c9;
         mem[1743] =  20'h010c9;
         mem[1744] =  20'h0a8d0;
         mem[1745] =  20'h068d0;
         mem[1746] =  20'h54cc9;
         mem[1747] =  20'h000c9;
         mem[1748] =  20'h218c6;
         mem[1749] =  20'h3f526;
         mem[1750] =  20'h2f470;
         mem[1751] =  20'h3f9cc;
         mem[1752] =  20'h27586;
         mem[1753] =  20'h0e494;
         mem[1754] =  20'h54cc9;
         mem[1755] =  20'h28089;
         mem[1756] =  20'h54cc9;
         mem[1757] =  20'h7e5c4;
         mem[1758] =  20'h1a20c;
         mem[1759] =  20'h27cc9;
         mem[1760] =  20'h00ea4;
         mem[1761] =  20'h524c9;
         mem[1762] =  20'h680a8;
         mem[1763] =  20'h01210;
         mem[1764] =  20'h271c6;
         mem[1765] =  20'h21c8f;
         mem[1766] =  20'h60188;
         mem[1767] =  20'h2d584;
         mem[1768] =  20'h26dc6;
         mem[1769] =  20'h2664a;
         mem[1770] =  20'h01a55;
         mem[1771] =  20'h00315;
         mem[1772] =  20'h72243;
         mem[1773] =  20'h5dd26;
         mem[1774] =  20'h13e62;
         mem[1775] =  20'h12f02;
         mem[1776] =  20'h5b524;
         mem[1777] =  20'h57924;
         mem[1778] =  20'h5f642;
         mem[1779] =  20'h6b243;
         mem[1780] =  20'h03077;
         mem[1781] =  20'h01906;
         mem[1782] =  20'h65a43;
         mem[1783] =  20'h02477;
         mem[1784] =  20'h2e48a;
         mem[1785] =  20'h33d4c;
         mem[1786] =  20'h3bcce;
         mem[1787] =  20'h00949;
         mem[1788] =  20'h090ac;
         mem[1789] =  20'h1958a;
         mem[1790] =  20'h0a124;
         mem[1791] =  20'h0cd0a;
         mem[1792] =  20'h08cac;
         mem[1793] =  20'h011d8;
         mem[1794] =  20'h6c144;
         mem[1795] =  20'h5a08a;
         mem[1796] =  20'h610c9;
         mem[1797] =  20'h84243;
         mem[1798] =  20'h610c9;
         mem[1799] =  20'h5f0c9;
         mem[1800] =  20'h28092;
         mem[1801] =  20'h148cb;
         mem[1802] =  20'h0a124;
         mem[1803] =  20'h1a5c8;
         mem[1804] =  20'h085e9;
         mem[1805] =  20'h0e50a;
         mem[1806] =  20'h0f8cc;
         mem[1807] =  20'h0e0cc;
         mem[1808] =  20'h2d984;
         mem[1809] =  20'h1458a;
         mem[1810] =  20'h26e06;
         mem[1811] =  20'h07249;
         mem[1812] =  20'h32e45;
         mem[1813] =  20'h00316;
         mem[1814] =  20'h67926;
         mem[1815] =  20'h64308;
         mem[1816] =  20'h772c4;
         mem[1817] =  20'h64526;
         mem[1818] =  20'h33d44;
         mem[1819] =  20'h600c9;
         mem[1820] =  20'h73186;
         mem[1821] =  20'h71186;
         mem[1822] =  20'h14e09;
         mem[1823] =  20'h1f546;
         mem[1824] =  20'h20a43;
         mem[1825] =  20'h26126;
         mem[1826] =  20'h10149;
         mem[1827] =  20'h26643;
         mem[1828] =  20'h0ede6;
         mem[1829] =  20'h331e6;
         mem[1830] =  20'h1f704;
         mem[1831] =  20'h33ccc;
         mem[1832] =  20'h02cc9;
         mem[1833] =  20'h4b0cc;
         mem[1834] =  20'h4e946;
         mem[1835] =  20'h2c649;
         mem[1836] =  20'h5a549;
         mem[1837] =  20'h27548;
         mem[1838] =  20'h271c6;
         mem[1839] =  20'h52527;
         mem[1840] =  20'h420cc;
         mem[1841] =  20'h3f8cc;
         mem[1842] =  20'h3b906;
         mem[1843] =  20'h14c8e;
         mem[1844] =  20'h04472;
         mem[1845] =  20'h4c20c;
         mem[1846] =  20'h03cce;
         mem[1847] =  20'h00cce;
         mem[1848] =  20'h0f994;
         mem[1849] =  20'h0c994;
         mem[1850] =  20'h040d1;
         mem[1851] =  20'h008d1;
         mem[1852] =  20'h29526;
         mem[1853] =  20'h25926;
         mem[1854] =  20'h0accd;
         mem[1855] =  20'h064cd;
         mem[1856] =  20'h04089;
         mem[1857] =  20'h3fd87;
         mem[1858] =  20'h3b586;
         mem[1859] =  20'h38586;
         mem[1860] =  20'h2d1c9;
         mem[1861] =  20'h5de83;
         mem[1862] =  20'h4090a;
         mem[1863] =  20'h1a5a9;
         mem[1864] =  20'h0f0d2;
         mem[1865] =  20'h018c9;
         mem[1866] =  20'h39d84;
         mem[1867] =  20'h0d5ec;
         mem[1868] =  20'h03185;
         mem[1869] =  20'h5de43;
         mem[1870] =  20'h57b05;
         mem[1871] =  20'h07872;
         mem[1872] =  20'h0288e;
         mem[1873] =  20'h15089;
         mem[1874] =  20'h0e986;
         mem[1875] =  20'h19224;
         mem[1876] =  20'h680a8;
         mem[1877] =  20'h64ca8;
         mem[1878] =  20'h72242;
         mem[1879] =  20'h00185;
         mem[1880] =  20'h164cc;
         mem[1881] =  20'h4b0cc;
         mem[1882] =  20'h136a3;
         mem[1883] =  20'h13ccc;
         mem[1884] =  20'h35186;
         mem[1885] =  20'h5de09;
         mem[1886] =  20'h52e45;
         mem[1887] =  20'h25de6;
         mem[1888] =  20'h3b126;
         mem[1889] =  20'h00deb;
         mem[1890] =  20'h16872;
         mem[1891] =  20'h14472;
         mem[1892] =  20'h21948;
         mem[1893] =  20'h1a208;
         mem[1894] =  20'h2d983;
         mem[1895] =  20'h0152d;
         mem[1896] =  20'h02cc9;
         mem[1897] =  20'h01cc9;
         mem[1898] =  20'h08549;
         mem[1899] =  20'h0ca42;
         mem[1900] =  20'h53dc6;
         mem[1901] =  20'h515c6;
         mem[1902] =  20'h11875;
         mem[1903] =  20'h384ac;
         mem[1904] =  20'h28986;
         mem[1905] =  20'h32683;
         mem[1906] =  20'h2d263;
         mem[1907] =  20'h4b526;
         mem[1908] =  20'h401cc;
         mem[1909] =  20'h26dd2;
         mem[1910] =  20'h4dd27;
         mem[1911] =  20'h5e244;
         mem[1912] =  20'h5a4c9;
         mem[1913] =  20'h32244;
         mem[1914] =  20'h3f686;
         mem[1915] =  20'h3ee86;
         mem[1916] =  20'h38702;
         mem[1917] =  20'h4b688;
         mem[1918] =  20'h4dd27;
         mem[1919] =  20'h4c127;
         mem[1920] =  20'h4e105;
         mem[1921] =  20'h4c105;
         mem[1922] =  20'h41c8a;
         mem[1923] =  20'h5e282;
         mem[1924] =  20'h40cc6;
         mem[1925] =  20'h066a3;
         mem[1926] =  20'h1a9a9;
         mem[1927] =  20'h20d85;
         mem[1928] =  20'h41146;
         mem[1929] =  20'h4c8a8;
         mem[1930] =  20'h034c9;
         mem[1931] =  20'h3f246;
         mem[1932] =  20'h0f524;
         mem[1933] =  20'h7d6a3;
         mem[1934] =  20'h3eec2;
         mem[1935] =  20'h6a643;
         mem[1936] =  20'h034c9;
         mem[1937] =  20'h014c9;
         mem[1938] =  20'h110d4;
         mem[1939] =  20'h0c8d4;
         mem[1940] =  20'h2e8ce;
         mem[1941] =  20'h06489;
         mem[1942] =  20'h5a924;
         mem[1943] =  20'h51924;
         mem[1944] =  20'h275e6;
         mem[1945] =  20'h0e872;
         mem[1946] =  20'h27186;
         mem[1947] =  20'h77684;
         mem[1948] =  20'h614c9;
         mem[1949] =  20'h2024e;
         mem[1950] =  20'h29492;
         mem[1951] =  20'h26c92;
         mem[1952] =  20'h02cc9;
         mem[1953] =  20'h01cc9;
         mem[1954] =  20'h220c9;
         mem[1955] =  20'h218c6;
         mem[1956] =  20'h07606;
         mem[1957] =  20'h538cb;
         mem[1958] =  20'h0a8cc;
         mem[1959] =  20'h6aa43;
         mem[1960] =  20'h53148;
         mem[1961] =  20'h72146;
         mem[1962] =  20'h59d24;
         mem[1963] =  20'h068cc;
         mem[1964] =  20'h1dcac;
         mem[1965] =  20'h00108;
         mem[1966] =  20'h20263;
         mem[1967] =  20'h1f986;
         mem[1968] =  20'h06ea8;
         mem[1969] =  20'h07608;
         mem[1970] =  20'h01a43;
         mem[1971] =  20'h1a14e;
         mem[1972] =  20'h2948a;
         mem[1973] =  20'h71643;
         mem[1974] =  20'h72986;
         mem[1975] =  20'h5e8c9;
         mem[1976] =  20'h2f8c8;
         mem[1977] =  20'h2c8c8;
         mem[1978] =  20'h39a46;
         mem[1979] =  20'h51986;
         mem[1980] =  20'h61546;
         mem[1981] =  20'h5dd46;
         mem[1982] =  20'h550c9;
         mem[1983] =  20'h520c9;
         mem[1984] =  20'h21908;
         mem[1985] =  20'h70d86;
         mem[1986] =  20'h7a144;
         mem[1987] =  20'h77144;
         mem[1988] =  20'h78643;
         mem[1989] =  20'h5988a;
         mem[1990] =  20'h00306;
         mem[1991] =  20'h064c9;
         mem[1992] =  20'h39686;
         mem[1993] =  20'h5e268;
         mem[1994] =  20'h03946;
         mem[1995] =  20'h3eeae;
         mem[1996] =  20'h41108;
         mem[1997] =  20'h33944;
         mem[1998] =  20'h21c89;
         mem[1999] =  20'h210ca;
         mem[2000] =  20'h1c88d;
         mem[2001] =  20'h1a88d;
         mem[2002] =  20'h2dd26;
         mem[2003] =  20'h26606;
         mem[2004] =  20'h1a60e;
         mem[2005] =  20'h00304;
         mem[2006] =  20'h08926;
         mem[2007] =  20'h075c4;
         mem[2008] =  20'h5a0e9;
         mem[2009] =  20'h14d0a;
         mem[2010] =  20'h14985;
         mem[2011] =  20'h0e88d;
         mem[2012] =  20'h0f473;
         mem[2013] =  20'h2d926;
         mem[2014] =  20'h8aa82;
         mem[2015] =  20'h64304;
         mem[2016] =  20'h14985;
         mem[2017] =  20'h3ed0e;
         mem[2018] =  20'h66cc6;
         mem[2019] =  20'h01958;
         mem[2020] =  20'h211ce;
         mem[2021] =  20'h33d48;
         mem[2022] =  20'h08926;
         mem[2023] =  20'h25b03;
         mem[2024] =  20'h14985;
         mem[2025] =  20'h51ac4;
         mem[2026] =  20'h4d586;
         mem[2027] =  20'h1f526;
         mem[2028] =  20'h1fae6;
         mem[2029] =  20'h25e6c;
         mem[2030] =  20'h088d5;
         mem[2031] =  20'h77a43;
         mem[2032] =  20'h59cc9;
         mem[2033] =  20'h27c8c;
         mem[2034] =  20'h040c9;
         mem[2035] =  20'h008c9;
         mem[2036] =  20'h09896;
         mem[2037] =  20'h3250c;
         mem[2038] =  20'h2f4e9;
         mem[2039] =  20'h4be44;
         mem[2040] =  20'h09896;
         mem[2041] =  20'h08096;
         mem[2042] =  20'h2ce84;
         mem[2043] =  20'h40cc7;
         mem[2044] =  20'h2d944;
         mem[2045] =  20'h12c8f;
         mem[2046] =  20'h03d0c;
         mem[2047] =  20'h0050c;
         mem[2048] =  20'h22cd0;
         mem[2049] =  20'h204d0;
         mem[2050] =  20'h03cd0;
         mem[2051] =  20'h00cd0;
         mem[2052] =  20'h0cb03;
         mem[2053] =  20'h08144;
         mem[2054] =  20'h006e8;
         mem[2055] =  20'h6aa63;
         mem[2056] =  20'h72242;
         mem[2057] =  20'h6a926;
         mem[2058] =  20'h618c9;
         mem[2059] =  20'h5e8c9;
         mem[2060] =  20'h58a86;
         mem[2061] =  20'h3e8ce;
         mem[2062] =  20'h72243;
         mem[2063] =  20'h4c127;
         mem[2064] =  20'h40245;
         mem[2065] =  20'h3ea45;
         mem[2066] =  20'h0d649;
         mem[2067] =  20'h2694a;
         mem[2068] =  20'h5c889;
         mem[2069] =  20'h57889;
         mem[2070] =  20'h09094;
         mem[2071] =  20'h84d83;
         mem[2072] =  20'h09094;
         mem[2073] =  20'h64548;
         mem[2074] =  20'h09094;
         mem[2075] =  20'h00473;
         mem[2076] =  20'h09094;
         mem[2077] =  20'h064c9;
         mem[2078] =  20'h2ca64;
         mem[2079] =  20'h59526;
         mem[2080] =  20'h0a8e6;
         mem[2081] =  20'h015c8;
         mem[2082] =  20'h0a506;
         mem[2083] =  20'h06506;
         mem[2084] =  20'h01a44;
         mem[2085] =  20'h57926;
         mem[2086] =  20'h2ca48;
         mem[2087] =  20'h454c9;
         mem[2088] =  20'h21cc9;
         mem[2089] =  20'h28092;
         mem[2090] =  20'h09094;
         mem[2091] =  20'h08894;
         mem[2092] =  20'h39a46;
         mem[2093] =  20'h1a8c9;
         mem[2094] =  20'h66906;
         mem[2095] =  20'h00248;
         mem[2096] =  20'h20dcc;
         mem[2097] =  20'h13de7;
         mem[2098] =  20'h4e946;
         mem[2099] =  20'h44c8a;
         mem[2100] =  20'h3eec3;
         mem[2101] =  20'h3a4ca;
         mem[2102] =  20'h0fccc;
         mem[2103] =  20'h28092;
         mem[2104] =  20'h33d50;
         mem[2105] =  20'h0850c;
         mem[2106] =  20'h0818e;
         mem[2107] =  20'h58186;
         mem[2108] =  20'h66cc6;
         mem[2109] =  20'h65cc6;
         mem[2110] =  20'h1c48a;
         mem[2111] =  20'h76e63;
         mem[2112] =  20'h350c8;
         mem[2113] =  20'h08516;
         mem[2114] =  20'h350c8;
         mem[2115] =  20'h338c8;
         mem[2116] =  20'h22cc9;
         mem[2117] =  20'h25b04;
         mem[2118] =  20'h4e946;
         mem[2119] =  20'h4b146;
         mem[2120] =  20'h26a63;
         mem[2121] =  20'h25e63;
         mem[2122] =  20'h01209;
         mem[2123] =  20'h06705;
         mem[2124] =  20'h264cf;
         mem[2125] =  20'h27cc9;
         mem[2126] =  20'h6a643;
         mem[2127] =  20'h8b242;
         mem[2128] =  20'h4b8c9;
         mem[2129] =  20'h4f8c9;
         mem[2130] =  20'h4b0c9;
         mem[2131] =  20'h5a48a;
         mem[2132] =  20'h27cd0;
         mem[2133] =  20'h2d94a;
         mem[2134] =  20'h130cd;
         mem[2135] =  20'h0accd;
         mem[2136] =  20'h078c9;
         mem[2137] =  20'h110cb;
         mem[2138] =  20'h0c8cb;
         mem[2139] =  20'h4d5e6;
         mem[2140] =  20'h0d283;
         mem[2141] =  20'h28089;
         mem[2142] =  20'h26d8e;
         mem[2143] =  20'h024c9;
         mem[2144] =  20'h01d26;
         mem[2145] =  20'h280c9;
         mem[2146] =  20'h07594;
         mem[2147] =  20'h2d643;
         mem[2148] =  20'h2be43;
         mem[2149] =  20'h7de43;
         mem[2150] =  20'h27cc9;
         mem[2151] =  20'h0e18f;
         mem[2152] =  20'h13643;
         mem[2153] =  20'h1dc92;
         mem[2154] =  20'h06663;
         mem[2155] =  20'h015e4;
         mem[2156] =  20'h0ddc5;
         mem[2157] =  20'h0cece;
         mem[2158] =  20'h5fcc9;
         mem[2159] =  20'h6be43;
         mem[2160] =  20'h27c72;
         mem[2161] =  20'h00a83;
         mem[2162] =  20'h1a4ac;
         mem[2163] =  20'h27985;
         mem[2164] =  20'h4d4cc;
         mem[2165] =  20'h5b10a;
         mem[2166] =  20'h5810a;
         mem[2167] =  20'h73186;
         mem[2168] =  20'h130c9;
         mem[2169] =  20'h15874;
         mem[2170] =  20'h269c6;
         mem[2171] =  20'h20d8d;
         mem[2172] =  20'h1a48f;
         mem[2173] =  20'h665e4;
         mem[2174] =  20'h33cce;
         mem[2175] =  20'h27546;
         mem[2176] =  20'h1fe43;
         mem[2177] =  20'h079e8;
         mem[2178] =  20'h08112;
         mem[2179] =  20'h3eb03;
         mem[2180] =  20'h0c8cd;
         mem[2181] =  20'h0410a;
         mem[2182] =  20'h07949;
         mem[2183] =  20'h26e43;
         mem[2184] =  20'h06703;
         mem[2185] =  20'h1bccb;
         mem[2186] =  20'h0010a;
         mem[2187] =  20'h65243;
         mem[2188] =  20'h64a43;
         mem[2189] =  20'h00e4a;
         mem[2190] =  20'h13695;
         mem[2191] =  20'h2d5c3;
         mem[2192] =  20'h38586;
         mem[2193] =  20'h586a4;
         mem[2194] =  20'h57aa4;
         mem[2195] =  20'h84a43;
         mem[2196] =  20'h83a43;
         mem[2197] =  20'h1dc92;
         mem[2198] =  20'h2ca43;
         mem[2199] =  20'h1dc92;
         mem[2200] =  20'h5f946;
         mem[2201] =  20'h53969;
         mem[2202] =  20'h2588a;
         mem[2203] =  20'h67d26;
         mem[2204] =  20'h1f892;
         mem[2205] =  20'h3450a;
         mem[2206] =  20'h33d0a;
         mem[2207] =  20'h34585;
         mem[2208] =  20'h33d27;
         mem[2209] =  20'h34585;
         mem[2210] =  20'h27527;
         mem[2211] =  20'h34585;
         mem[2212] =  20'h21c92;
         mem[2213] =  20'h209cc;
         mem[2214] =  20'h06564;
         mem[2215] =  20'h40cca;
         mem[2216] =  20'h6ad66;
         mem[2217] =  20'h67d26;
         mem[2218] =  20'h3ee42;
         mem[2219] =  20'h1a98d;
         mem[2220] =  20'h70a43;
         mem[2221] =  20'h72243;
         mem[2222] =  20'h64126;
         mem[2223] =  20'h61126;
         mem[2224] =  20'h5e526;
         mem[2225] =  20'h098d0;
         mem[2226] =  20'h078d0;
         mem[2227] =  20'h220ca;
         mem[2228] =  20'h210ca;
         mem[2229] =  20'h028d8;
         mem[2230] =  20'h19c94;
         mem[2231] =  20'h038c9;
         mem[2232] =  20'h010c9;
         mem[2233] =  20'h20645;
         mem[2234] =  20'h26cc9;
         mem[2235] =  20'h0e5e8;
         mem[2236] =  20'h0d1e8;
         mem[2237] =  20'h02889;
         mem[2238] =  20'h19ccc;
         mem[2239] =  20'h04112;
         mem[2240] =  20'h00112;
         mem[2241] =  20'h2bf06;
         mem[2242] =  20'h2cdc3;
         mem[2243] =  20'h3490f;
         mem[2244] =  20'h01d4e;
         mem[2245] =  20'h41d0a;
         mem[2246] =  20'h00c89;
         mem[2247] =  20'h0a4c8;
         mem[2248] =  20'h06cc8;
         mem[2249] =  20'h2664c;
         mem[2250] =  20'h4c204;
         mem[2251] =  20'h3960f;
         mem[2252] =  20'h3f50a;
         mem[2253] =  20'h72a06;
         mem[2254] =  20'h64985;
         mem[2255] =  20'h5b124;
         mem[2256] =  20'h59526;
         mem[2257] =  20'h3fa0c;
         mem[2258] =  20'h51666;
         mem[2259] =  20'h53d26;
         mem[2260] =  20'h01477;
         mem[2261] =  20'h32306;
         mem[2262] =  20'h1f4ac;
         mem[2263] =  20'h00e72;
         mem[2264] =  20'h470cc;
         mem[2265] =  20'h1f708;
         mem[2266] =  20'h72124;
         mem[2267] =  20'h34146;
         mem[2268] =  20'h2c683;
         mem[2269] =  20'h030f4;
         mem[2270] =  20'h014f4;
         mem[2271] =  20'h10052;
         mem[2272] =  20'h3354c;
         mem[2273] =  20'h39d88;
         mem[2274] =  20'h2d86e;
         mem[2275] =  20'h0f590;
         mem[2276] =  20'h01cc9;
         mem[2277] =  20'h5ad24;
         mem[2278] =  20'h4b2c4;
         mem[2279] =  20'h4b6c6;
         mem[2280] =  20'h27126;
         mem[2281] =  20'h02889;
         mem[2282] =  20'h32e47;
         mem[2283] =  20'h25b06;
         mem[2284] =  20'h44f0a;
         mem[2285] =  20'h13a55;
         mem[2286] =  20'h4cc8a;
         mem[2287] =  20'h66948;
         mem[2288] =  20'h278c9;
         mem[2289] =  20'h418cc;
         mem[2290] =  20'h400cc;
         mem[2291] =  20'h4f0cc;
         mem[2292] =  20'h4b8cc;
         mem[2293] =  20'h604c9;
         mem[2294] =  20'h5fcc9;
         mem[2295] =  20'h80944;
         mem[2296] =  20'h7d144;
         mem[2297] =  20'h6d126;
         mem[2298] =  20'h0d5c4;
         mem[2299] =  20'h08d44;
         mem[2300] =  20'h5dd44;
         mem[2301] =  20'h11473;
         mem[2302] =  20'h4c128;
         mem[2303] =  20'h2ccac;
         mem[2304] =  20'h06703;
         mem[2305] =  20'h33984;
         mem[2306] =  20'h1788a;
         mem[2307] =  20'h25926;
         mem[2308] =  20'h048d6;
         mem[2309] =  20'h000d6;
         mem[2310] =  20'h5f263;
         mem[2311] =  20'h2e48f;
         mem[2312] =  20'h27cc9;
         mem[2313] =  20'h83643;
         mem[2314] =  20'h1494f;
         mem[2315] =  20'h2c243;
         mem[2316] =  20'h0e926;
         mem[2317] =  20'h3eb0e;
         mem[2318] =  20'h3b90a;
         mem[2319] =  20'h21c89;
         mem[2320] =  20'h3b90a;
         mem[2321] =  20'h4694a;
         mem[2322] =  20'h52644;
         mem[2323] =  20'h00262;
         mem[2324] =  20'h70b06;
         mem[2325] =  20'h1a910;
         mem[2326] =  20'h33d44;
         mem[2327] =  20'h12cc9;
         mem[2328] =  20'h610e9;
         mem[2329] =  20'h71586;
         mem[2330] =  20'h5a8c9;
         mem[2331] =  20'h5e5e8;
         mem[2332] =  20'h27cd0;
         mem[2333] =  20'h270ec;
         mem[2334] =  20'h290c9;
         mem[2335] =  20'h58cc9;
         mem[2336] =  20'h348c9;
         mem[2337] =  20'h27092;
         mem[2338] =  20'h3bccc;
         mem[2339] =  20'h394cc;
         mem[2340] =  20'h61526;
         mem[2341] =  20'h7d244;
         mem[2342] =  20'h73d26;
         mem[2343] =  20'h71126;
         mem[2344] =  20'h65a43;
         mem[2345] =  20'h64243;
         mem[2346] =  20'h11496;
         mem[2347] =  20'h0cc96;
         mem[2348] =  20'h03c58;
         mem[2349] =  20'h7de04;
         mem[2350] =  20'h28492;
         mem[2351] =  20'h3a14e;
         mem[2352] =  20'h290c9;
         mem[2353] =  20'h264e9;
         mem[2354] =  20'h1e094;
         mem[2355] =  20'h274c9;
         mem[2356] =  20'h01d4e;
         mem[2357] =  20'h06e46;
         mem[2358] =  20'h03c58;
         mem[2359] =  20'h01c58;
         mem[2360] =  20'h4e4c7;
         mem[2361] =  20'h4c4c7;
         mem[2362] =  20'h20253;
         mem[2363] =  20'h26d26;
         mem[2364] =  20'h21926;
         mem[2365] =  20'h64d48;
         mem[2366] =  20'h36caf;
         mem[2367] =  20'h320af;
         mem[2368] =  20'h1e094;
         mem[2369] =  20'h19094;
         mem[2370] =  20'h2d944;
         mem[2371] =  20'h77dc4;
         mem[2372] =  20'h47583;
         mem[2373] =  20'h06703;
         mem[2374] =  20'h0e5d4;
         mem[2375] =  20'h514c9;
         mem[2376] =  20'h03493;
         mem[2377] =  20'h451c3;
         mem[2378] =  20'h08214;
         mem[2379] =  20'h3eaa9;
         mem[2380] =  20'h785e5;
         mem[2381] =  20'h408c6;
         mem[2382] =  20'h08214;
         mem[2383] =  20'h06a14;
         mem[2384] =  20'h1d06c;
         mem[2385] =  20'h1a46c;
         mem[2386] =  20'h27548;
         mem[2387] =  20'h394c6;
         mem[2388] =  20'h20d84;
         mem[2389] =  20'h0ecaf;
         mem[2390] =  20'h03d26;
         mem[2391] =  20'h0196a;
         mem[2392] =  20'h2ec8c;
         mem[2393] =  20'h0e524;
         mem[2394] =  20'h019a6;
         mem[2395] =  20'h28092;
         mem[2396] =  20'h348c9;
         mem[2397] =  20'h71546;
         mem[2398] =  20'h58a83;
         mem[2399] =  20'h5e526;
         mem[2400] =  20'h03493;
         mem[2401] =  20'h01c93;
         mem[2402] =  20'h196c2;
         mem[2403] =  20'h00126;
         mem[2404] =  20'h00312;
         mem[2405] =  20'h0d608;
         mem[2406] =  20'h26646;
         mem[2407] =  20'h070ca;
         mem[2408] =  20'h03526;
         mem[2409] =  20'h00926;
         mem[2410] =  20'h0f08f;
         mem[2411] =  20'h018ea;
         mem[2412] =  20'h0d284;
         mem[2413] =  20'h45663;
         mem[2414] =  20'h348c9;
         mem[2415] =  20'h340c9;
         mem[2416] =  20'h35489;
         mem[2417] =  20'h45929;
         mem[2418] =  20'h39245;
         mem[2419] =  20'h19854;
         mem[2420] =  20'h6dd06;
         mem[2421] =  20'h84242;
         mem[2422] =  20'h1a5e6;
         mem[2423] =  20'h5e586;
         mem[2424] =  20'h364c9;
         mem[2425] =  20'h4ba84;
         mem[2426] =  20'h6a706;
         mem[2427] =  20'h65d24;
         mem[2428] =  20'h0a096;
         mem[2429] =  20'h07896;
         mem[2430] =  20'h54109;
         mem[2431] =  20'h07cc9;
         mem[2432] =  20'h1bc72;
         mem[2433] =  20'h33586;
         mem[2434] =  20'h2f8a8;
         mem[2435] =  20'h2cca8;
         mem[2436] =  20'h288cc;
         mem[2437] =  20'h270cc;
         mem[2438] =  20'h399c8;
         mem[2439] =  20'h0886e;
         mem[2440] =  20'h288cc;
         mem[2441] =  20'h20492;
         mem[2442] =  20'h26a12;
         mem[2443] =  20'h1a4f4;
         mem[2444] =  20'h3590c;
         mem[2445] =  20'h40cce;
         mem[2446] =  20'h21926;
         mem[2447] =  20'h1b472;
         mem[2448] =  20'h196ce;
         mem[2449] =  20'h2c642;
         mem[2450] =  20'h288cc;
         mem[2451] =  20'h20d27;
         mem[2452] =  20'h2ec8c;
         mem[2453] =  20'h2dc8c;
         mem[2454] =  20'h0e556;
         mem[2455] =  20'h06474;
         mem[2456] =  20'h52644;
         mem[2457] =  20'h51e44;
         mem[2458] =  20'h61926;
         mem[2459] =  20'h5dd26;
         mem[2460] =  20'h01a58;
         mem[2461] =  20'h270cc;
         mem[2462] =  20'h2dd44;
         mem[2463] =  20'h38a46;
         mem[2464] =  20'h27243;
         mem[2465] =  20'h2d928;
         mem[2466] =  20'h4d8cc;
         mem[2467] =  20'h58643;
         mem[2468] =  20'h6e127;
         mem[2469] =  20'h4b546;
         mem[2470] =  20'h6e127;
         mem[2471] =  20'h15473;
         mem[2472] =  20'h6e127;
         mem[2473] =  20'h07d69;
         mem[2474] =  20'h6e127;
         mem[2475] =  20'h20d66;
         mem[2476] =  20'h2fd05;
         mem[2477] =  20'h19a93;
         mem[2478] =  20'h06ea6;
         mem[2479] =  20'h20d8e;
         mem[2480] =  20'h024c9;
         mem[2481] =  20'h45505;
         mem[2482] =  20'h2fd05;
         mem[2483] =  20'h2bd05;
         mem[2484] =  20'h6e127;
         mem[2485] =  20'h2790a;
         mem[2486] =  20'h61929;
         mem[2487] =  20'h5dd29;
         mem[2488] =  20'h41927;
         mem[2489] =  20'h3f527;
         mem[2490] =  20'h61148;
         mem[2491] =  20'h064cc;
         mem[2492] =  20'h028cc;
         mem[2493] =  20'h01d4c;
         mem[2494] =  20'h07608;
         mem[2495] =  20'h83663;
         mem[2496] =  20'h39e44;
         mem[2497] =  20'h19d26;
         mem[2498] =  20'h088cf;
         mem[2499] =  20'h398c6;
         mem[2500] =  20'h079c9;
         mem[2501] =  20'h00d14;
         mem[2502] =  20'h014e9;
         mem[2503] =  20'h27185;
         mem[2504] =  20'h0650e;
         mem[2505] =  20'h4bac4;
         mem[2506] =  20'h6c4c6;
         mem[2507] =  20'h0acc7;
         mem[2508] =  20'h000c6;
         mem[2509] =  20'h26a32;
         mem[2510] =  20'h01986;
         mem[2511] =  20'h2ce44;
         mem[2512] =  20'h4c146;
         mem[2513] =  20'h3a14c;
         mem[2514] =  20'h06703;
         mem[2515] =  20'h480c6;
         mem[2516] =  20'h460c6;
         mem[2517] =  20'h3f663;
         mem[2518] =  20'h0c8c9;
         mem[2519] =  20'h67946;
         mem[2520] =  20'h64146;
         mem[2521] =  20'h54d26;
         mem[2522] =  20'h64243;
         mem[2523] =  20'h65a43;
         mem[2524] =  20'h70926;
         mem[2525] =  20'h54d26;
         mem[2526] =  20'h0e0c9;
         mem[2527] =  20'h35c8c;
         mem[2528] =  20'h53508;
         mem[2529] =  20'h7e243;
         mem[2530] =  20'h3348c;
         mem[2531] =  20'h2d983;
         mem[2532] =  20'h28089;
         mem[2533] =  20'h7e643;
         mem[2534] =  20'h7d643;
         mem[2535] =  20'h0acd4;
         mem[2536] =  20'h064d4;
         mem[2537] =  20'h16092;
         mem[2538] =  20'h0c8cc;
         mem[2539] =  20'h3b586;
         mem[2540] =  20'h14892;
         mem[2541] =  20'h038c9;
         mem[2542] =  20'h38586;
         mem[2543] =  20'h1c914;
         mem[2544] =  20'h19914;
         mem[2545] =  20'h54d26;
         mem[2546] =  20'h51926;
         mem[2547] =  20'h5ea43;
         mem[2548] =  20'h52926;
         mem[2549] =  20'h01643;
         mem[2550] =  20'h0e8c7;
         mem[2551] =  20'h08926;
         mem[2552] =  20'h07d26;
         mem[2553] =  20'h26dc6;
         mem[2554] =  20'h0e8cd;
         mem[2555] =  20'h46586;
         mem[2556] =  20'h0724f;
         mem[2557] =  20'h034c7;
         mem[2558] =  20'h13a06;
         mem[2559] =  20'h0946c;
         mem[2560] =  20'h2d8c9;
         mem[2561] =  20'h03498;
         mem[2562] =  20'h01c98;
         mem[2563] =  20'h3b0ac;
         mem[2564] =  20'h5f926;
         mem[2565] =  20'h2d246;
         mem[2566] =  20'h3a4ac;
         mem[2567] =  20'h6b626;
         mem[2568] =  20'h12e4e;
         mem[2569] =  20'h06702;
         mem[2570] =  20'h5de43;
         mem[2571] =  20'h024c9;
         mem[2572] =  20'h139cc;
         mem[2573] =  20'h0946c;
         mem[2574] =  20'h020c9;
         mem[2575] =  20'h280ca;
         mem[2576] =  20'h014c9;
         mem[2577] =  20'h00aa7;
         mem[2578] =  20'h46585;
         mem[2579] =  20'h2dd28;
         mem[2580] =  20'h27cd2;
         mem[2581] =  20'h5b50a;
         mem[2582] =  20'h57d0a;
         mem[2583] =  20'h02d0a;
         mem[2584] =  20'h0150a;
         mem[2585] =  20'h07d85;
         mem[2586] =  20'h4b642;
         mem[2587] =  20'h32a86;
         mem[2588] =  20'h27527;
         mem[2589] =  20'h21d10;
         mem[2590] =  20'h39208;
         mem[2591] =  20'h33d44;
         mem[2592] =  20'h4cd48;
         mem[2593] =  20'h791e4;
         mem[2594] =  20'h00649;
         mem[2595] =  20'h1c548;
         mem[2596] =  20'h64e44;
         mem[2597] =  20'h2dd4c;
         mem[2598] =  20'h2d54c;
         mem[2599] =  20'h26a47;
         mem[2600] =  20'h6a643;
         mem[2601] =  20'h6b243;
         mem[2602] =  20'h198ca;
         mem[2603] =  20'h04118;
         mem[2604] =  20'h0110f;
         mem[2605] =  20'h04118;
         mem[2606] =  20'h19649;
         mem[2607] =  20'h4ed26;
         mem[2608] =  20'h39246;
         mem[2609] =  20'h23cc9;
         mem[2610] =  20'h1f4c9;
         mem[2611] =  20'h2ce44;
         mem[2612] =  20'h06d94;
         mem[2613] =  20'h044d7;
         mem[2614] =  20'h25c52;
         mem[2615] =  20'h34146;
         mem[2616] =  20'h25a86;
         mem[2617] =  20'h4dd85;
         mem[2618] =  20'h19073;
         mem[2619] =  20'h0b072;
         mem[2620] =  20'h06c72;
         mem[2621] =  20'h3f643;
         mem[2622] =  20'h1a149;
         mem[2623] =  20'h531c7;
         mem[2624] =  20'h521c7;
         mem[2625] =  20'h5fd26;
         mem[2626] =  20'h5890a;
         mem[2627] =  20'h5a08a;
         mem[2628] =  20'h32cb0;
         mem[2629] =  20'h42526;
         mem[2630] =  20'h3e926;
         mem[2631] =  20'h2d589;
         mem[2632] =  20'h40ca8;
         mem[2633] =  20'h0946c;
         mem[2634] =  20'h5fcc9;
         mem[2635] =  20'h298e6;
         mem[2636] =  20'h08496;
         mem[2637] =  20'h271c3;
         mem[2638] =  20'h70a63;
         mem[2639] =  20'h044d8;
         mem[2640] =  20'h515e6;
         mem[2641] =  20'h27d4e;
         mem[2642] =  20'h25d0a;
         mem[2643] =  20'h27585;
         mem[2644] =  20'h2d926;
         mem[2645] =  20'h33dce;
         mem[2646] =  20'h32dce;
         mem[2647] =  20'h345a4;
         mem[2648] =  20'h0d4cc;
         mem[2649] =  20'h40226;
         mem[2650] =  20'h3ee26;
         mem[2651] =  20'h2fd09;
         mem[2652] =  20'h2bd09;
         mem[2653] =  20'h3870a;
         mem[2654] =  20'h0d5e8;
         mem[2655] =  20'h0da48;
         mem[2656] =  20'h06644;
         mem[2657] =  20'h11872;
         mem[2658] =  20'h13073;
         mem[2659] =  20'h368d0;
         mem[2660] =  20'h320d0;
         mem[2661] =  20'h72966;
         mem[2662] =  20'h26985;
         mem[2663] =  20'h27585;
         mem[2664] =  20'h14526;
         mem[2665] =  20'h27585;
         mem[2666] =  20'h344c7;
         mem[2667] =  20'h0e926;
         mem[2668] =  20'h598c9;
         mem[2669] =  20'h0e926;
         mem[2670] =  20'h13e14;
         mem[2671] =  20'h2754c;
         mem[2672] =  20'h0c8ec;
         mem[2673] =  20'h6d566;
         mem[2674] =  20'h2cd88;
         mem[2675] =  20'h46d0a;
         mem[2676] =  20'h08889;
         mem[2677] =  20'h03876;
         mem[2678] =  20'h01c76;
         mem[2679] =  20'h2ce44;
         mem[2680] =  20'h0f08f;
         mem[2681] =  20'h0946c;
         mem[2682] =  20'h0024d;
         mem[2683] =  20'h04078;
         mem[2684] =  20'h01478;
         mem[2685] =  20'h604a8;
         mem[2686] =  20'h71242;
         mem[2687] =  20'h32a83;
         mem[2688] =  20'h27526;
         mem[2689] =  20'h0d66a;
         mem[2690] =  20'h2c663;
         mem[2691] =  20'h29524;
         mem[2692] =  20'h0d248;
         mem[2693] =  20'h3adc4;
         mem[2694] =  20'h1a0d0;
         mem[2695] =  20'h35d30;
         mem[2696] =  20'h32130;
         mem[2697] =  20'h048ce;
         mem[2698] =  20'h000ce;
         mem[2699] =  20'h03cd6;
         mem[2700] =  20'h00cd6;
         mem[2701] =  20'h0f994;
         mem[2702] =  20'h0c994;
         mem[2703] =  20'h28489;
         mem[2704] =  20'h024d0;
         mem[2705] =  20'h0946c;
         mem[2706] =  20'h19e46;
         mem[2707] =  20'h20a08;
         mem[2708] =  20'h51546;
         mem[2709] =  20'h59926;
         mem[2710] =  20'h0e126;
         mem[2711] =  20'h09d48;
         mem[2712] =  20'h0886c;
         mem[2713] =  20'h1a989;
         mem[2714] =  20'h20d86;
         mem[2715] =  20'h06905;
         mem[2716] =  20'h4e0c8;
         mem[2717] =  20'h4bd86;
         mem[2718] =  20'h72d86;
         mem[2719] =  20'h524c6;
         mem[2720] =  20'h158f2;
         mem[2721] =  20'h39243;
         mem[2722] =  20'h14262;
         mem[2723] =  20'h0d986;
         mem[2724] =  20'h27cc9;
         mem[2725] =  20'h278c9;
         mem[2726] =  20'h3c4af;
         mem[2727] =  20'h390af;
         mem[2728] =  20'h271c6;
         mem[2729] =  20'h2786e;
         mem[2730] =  20'h64305;
         mem[2731] =  20'h7d283;
         mem[2732] =  20'h3fe42;
         mem[2733] =  20'h258ca;
         mem[2734] =  20'h06e83;
         mem[2735] =  20'h538cb;
         mem[2736] =  20'h600c8;
         mem[2737] =  20'h4d4c9;
         mem[2738] =  20'h46242;
         mem[2739] =  20'h261e6;
         mem[2740] =  20'h01a43;
         mem[2741] =  20'h01472;
         mem[2742] =  20'h174ca;
         mem[2743] =  20'h12cca;
         mem[2744] =  20'h21d09;
         mem[2745] =  20'h20d09;
         mem[2746] =  20'h0d683;
         mem[2747] =  20'h0dda4;
         mem[2748] =  20'h044ee;
         mem[2749] =  20'h000ee;
         mem[2750] =  20'h47146;
         mem[2751] =  20'h46146;
         mem[2752] =  20'h28472;
         mem[2753] =  20'h64243;
         mem[2754] =  20'h65a43;
         mem[2755] =  20'h2692a;
         mem[2756] =  20'h2e1e4;
         mem[2757] =  20'h26d86;
         mem[2758] =  20'h07d89;
         mem[2759] =  20'h3a0cc;
         mem[2760] =  20'h221a6;
         mem[2761] =  20'h452cd;
         mem[2762] =  20'h368c6;
         mem[2763] =  20'h320c6;
         mem[2764] =  20'h25b03;
         mem[2765] =  20'h1f546;
         mem[2766] =  20'h2d643;
         mem[2767] =  20'h00146;
         mem[2768] =  20'h04c73;
         mem[2769] =  20'h26990;
         mem[2770] =  20'h2a492;
         mem[2771] =  20'h25c92;
         mem[2772] =  20'h84243;
         mem[2773] =  20'h76d24;
         mem[2774] =  20'h73986;
         mem[2775] =  20'h72524;
         mem[2776] =  20'h67148;
         mem[2777] =  20'h64948;
         mem[2778] =  20'h0394c;
         mem[2779] =  20'h0014c;
         mem[2780] =  20'h5b526;
         mem[2781] =  20'h57926;
         mem[2782] =  20'h5b146;
         mem[2783] =  20'h57946;
         mem[2784] =  20'h71e42;
         mem[2785] =  20'h70a43;
         mem[2786] =  20'h2024c;
         mem[2787] =  20'h140e9;
         mem[2788] =  20'h0126f;
         mem[2789] =  20'h00e04;
         mem[2790] =  20'h4c20c;
         mem[2791] =  20'h13d8f;
         mem[2792] =  20'h1d053;
         mem[2793] =  20'h1a853;
         mem[2794] =  20'h5ad0a;
         mem[2795] =  20'h5850a;
         mem[2796] =  20'h28872;
         mem[2797] =  20'h46186;
         mem[2798] =  20'h21d0a;
         mem[2799] =  20'h1a98a;
         mem[2800] =  20'h33a4a;
         mem[2801] =  20'h3224a;
         mem[2802] =  20'h28872;
         mem[2803] =  20'h57a43;
         mem[2804] =  20'h28872;
         mem[2805] =  20'h27c72;
         mem[2806] =  20'h59243;
         mem[2807] =  20'h1f643;
         mem[2808] =  20'h1fec3;
         mem[2809] =  20'h002aa;
         mem[2810] =  20'h14651;
         mem[2811] =  20'h12e51;
         mem[2812] =  20'h4b30b;
         mem[2813] =  20'h3fa06;
         mem[2814] =  20'h350c8;
         mem[2815] =  20'h59107;
         mem[2816] =  20'h424ce;
         mem[2817] =  20'h3f4ce;
         mem[2818] =  20'h4ca42;
         mem[2819] =  20'h33546;
         mem[2820] =  20'h47d24;
         mem[2821] =  20'h44d26;
         mem[2822] =  20'h0f472;
         mem[2823] =  20'h0f072;
         mem[2824] =  20'h4d4ca;
         mem[2825] =  20'h3ecc9;
         mem[2826] =  20'h39e06;
         mem[2827] =  20'h32526;
         mem[2828] =  20'h2da06;
         mem[2829] =  20'h00243;
         mem[2830] =  20'h028c9;
         mem[2831] =  20'h218c6;
         mem[2832] =  20'h28092;
         mem[2833] =  20'h020c9;
         mem[2834] =  20'h088c9;
         mem[2835] =  20'h00649;
         mem[2836] =  20'h12f03;
         mem[2837] =  20'h59124;
         mem[2838] =  20'h3a50a;
         mem[2839] =  20'h0dda9;
         mem[2840] =  20'h1a209;
         mem[2841] =  20'h1a1c9;
         mem[2842] =  20'h21526;
         mem[2843] =  20'h2c206;
         mem[2844] =  20'h21da9;
         mem[2845] =  20'h1f9a9;
         mem[2846] =  20'h19306;
         mem[2847] =  20'h57d49;
         mem[2848] =  20'h6ba43;
         mem[2849] =  20'h64243;
         mem[2850] =  20'h6c926;
         mem[2851] =  20'h7d6c4;
         mem[2852] =  20'h59906;
         mem[2853] =  20'h2790f;
         mem[2854] =  20'h1a643;
         mem[2855] =  20'h150aa;
         mem[2856] =  20'h33983;
         mem[2857] =  20'h26246;
         mem[2858] =  20'h28092;
         mem[2859] =  20'h210c6;
         mem[2860] =  20'h22c52;
         mem[2861] =  20'h21452;
         mem[2862] =  20'h0ed46;
         mem[2863] =  20'h0724c;
         mem[2864] =  20'h0de36;
         mem[2865] =  20'h01186;
         mem[2866] =  20'h39e06;
         mem[2867] =  20'h024b2;
         mem[2868] =  20'h030c9;
         mem[2869] =  20'h018c9;
         mem[2870] =  20'h088cc;
         mem[2871] =  20'h399a4;
         mem[2872] =  20'h33663;
         mem[2873] =  20'h3a8c8;
         mem[2874] =  20'h3b08f;
         mem[2875] =  20'h008ce;
         mem[2876] =  20'h0a0ce;
         mem[2877] =  20'h070ce;
         mem[2878] =  20'h7de44;
         mem[2879] =  20'h01494;
         mem[2880] =  20'h3610c;
         mem[2881] =  20'h3210c;
         mem[2882] =  20'h54948;
         mem[2883] =  20'h51948;
         mem[2884] =  20'h35c8f;
         mem[2885] =  20'h3348f;
         mem[2886] =  20'h4660c;
         mem[2887] =  20'h4560c;
         mem[2888] =  20'h4e8e9;
         mem[2889] =  20'h08c75;
         mem[2890] =  20'h48124;
         mem[2891] =  20'h3f629;
         mem[2892] =  20'h3550f;
         mem[2893] =  20'h32d0f;
         mem[2894] =  20'h5a548;
         mem[2895] =  20'h70ac6;
         mem[2896] =  20'h64304;
         mem[2897] =  20'h7e983;
         mem[2898] =  20'h4f8cc;
         mem[2899] =  20'h4b0cc;
         mem[2900] =  20'h6e126;
         mem[2901] =  20'h25eca;
         mem[2902] =  20'h6e126;
         mem[2903] =  20'h70a42;
         mem[2904] =  20'h5ea63;
         mem[2905] =  20'h51643;
         mem[2906] =  20'h6e126;
         mem[2907] =  20'h6a526;
         mem[2908] =  20'h6d526;
         mem[2909] =  20'h6b126;
         mem[2910] =  20'h10874;
         mem[2911] =  20'h51708;
         mem[2912] =  20'h088d6;
     end

endmodule: rect0_rom
